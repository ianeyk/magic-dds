magic
tech sky130A
timestamp 1702371875
<< locali >>
rect -130 7810 0 7830
rect -130 6655 -110 7810
rect -150 6635 -110 6655
rect -40 6520 0 6530
rect -40 6500 -30 6520
rect -10 6500 0 6520
rect -40 6490 0 6500
rect -150 5330 -95 5340
rect -150 5320 -125 5330
rect -135 5310 -125 5320
rect -105 5310 -95 5330
rect -135 5300 -95 5310
rect -135 5190 0 5200
rect -135 5170 -125 5190
rect -105 5180 0 5190
rect -105 5170 -95 5180
rect -135 5160 -95 5170
rect -150 4005 -110 4025
rect -130 3885 -110 4005
rect -130 3865 0 3885
rect -135 2720 -95 2730
rect -135 2710 -125 2720
rect -150 2700 -125 2710
rect -105 2700 -95 2720
rect -150 2690 -95 2700
rect -95 2580 -55 2590
rect -95 2560 -85 2580
rect -65 2570 -55 2580
rect -65 2560 0 2570
rect -95 2550 0 2560
rect -65 1405 -25 1415
rect -65 1395 -55 1405
rect -150 1385 -55 1395
rect -35 1385 -25 1405
rect -150 1375 -25 1385
rect -130 1235 0 1255
rect -130 80 -110 1235
rect -150 60 -110 80
<< viali >>
rect -30 6500 -10 6520
rect -125 5310 -105 5330
rect -125 5170 -105 5190
rect -125 2700 -105 2720
rect -85 2560 -65 2580
rect -55 1385 -35 1405
<< metal1 >>
rect -40 6520 0 6530
rect -40 6500 -30 6520
rect -10 6500 0 6520
rect -40 6490 0 6500
rect -135 5330 -95 5340
rect -135 5310 -125 5330
rect -105 5315 -95 5330
rect -105 5310 -65 5315
rect -135 5300 -65 5310
rect -135 5190 -95 5200
rect -135 5170 -125 5190
rect -105 5170 -95 5190
rect -135 5160 -95 5170
rect -135 2730 -120 5160
rect -135 2720 -95 2730
rect -135 2700 -125 2720
rect -105 2700 -95 2720
rect -135 2690 -95 2700
rect -80 2590 -65 5300
rect -95 2580 -55 2590
rect -95 2560 -85 2580
rect -65 2560 -55 2580
rect -95 2550 -55 2560
rect -40 1415 -25 6490
rect -65 1405 -25 1415
rect -65 1385 -55 1405
rect -35 1385 -25 1405
rect -65 1375 -25 1385
use half_dac_for_mirroring  half_dac_for_mirroring_0
timestamp 1702367632
transform 1 0 650 0 1 1315
box -650 -1315 2600 6575
use half_dac_for_mirroring  half_dac_for_mirroring_1
timestamp 1702367632
transform -1 0 -800 0 -1 6575
box -650 -1315 2600 6575
<< end >>
