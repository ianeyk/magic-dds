* SPICE3 file created from current_steering_dac.ext - technology: sky130A

.subckt dummy_current_steering_dac_unit_cell_with_encoder I1 I2 Vbn Vcn Vx Vx1 Vy
+ VP VN VN2
X0 a_200_0# Vbn VN2 VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X1 a_870_2050# Vy VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X2 a_530_1630# Vy a_560_2180# VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X3 VP Vx a_870_2050# VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 a_400_0# Vcn a_200_0# VN sky130_fd_pr__nfet_01v8 ad=3.3 pd=12.7 as=3 ps=12.5 w=12 l=0.5
X5 VP a_530_1630# a_560_1530# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X6 a_560_2180# Vx VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X7 a_870_2050# Vx1 a_530_1630# VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X8 VN a_530_1630# a_560_1530# VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X9 I1 VN a_400_0# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=2.2 ps=8.46 w=3 l=0.5
X10 VN Vx1 a_530_1630# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X11 I2 VN a_400_0# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=2.2 ps=8.46 w=3 l=0.5
.ends

.subckt current_steering_dac_unit_cell_with_encoder I1 I2 Vbn Vcn Vx Vx1 Vy VP VN
+ VN2
X0 a_200_0# Vbn VN2 VN sky130_fd_pr__nfet_01v8 ad=3 pd=12.5 as=6 ps=25 w=12 l=0.5
X1 a_870_2050# Vy VP VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X2 a_520_760# Vy a_560_2180# VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X3 VP Vx a_870_2050# VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X4 a_400_0# Vcn a_200_0# VN sky130_fd_pr__nfet_01v8 ad=2.2 pd=8.46 as=3 ps=12.5 w=12 l=0.5
X5 VP a_520_760# a_520_n30# VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X6 a_560_2180# Vx VN VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X7 a_870_2050# Vx1 a_520_760# VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X8 VN a_520_760# a_520_n30# VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.5 ps=3 w=1 l=0.15
X9 I1 a_520_n30# a_400_0# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=2.2 ps=8.46 w=3 l=0.5
X10 VN Vx1 a_520_760# VN sky130_fd_pr__nfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X11 I2 a_520_760# a_400_0# VN sky130_fd_pr__nfet_01v8 ad=1.5 pd=7 as=2.2 ps=8.46 w=3 l=0.5
.ends

.subckt half_dac_for_mirroring dummy_current_steering_dac_unit_cell_with_encoder_4/Vx1
+ current_steering_dac_unit_cell_with_encoder_6/VN2 dummy_current_steering_dac_unit_cell_with_encoder_1/Vx1
+ current_steering_dac_unit_cell_with_encoder_6/Vx1 current_steering_dac_unit_cell_with_encoder_8/Vbn
+ current_steering_dac_unit_cell_with_encoder_8/Vcn dummy_current_steering_dac_unit_cell_with_encoder_2/Vx1
+ current_steering_dac_unit_cell_with_encoder_9/VP current_steering_dac_unit_cell_with_encoder_8/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder_13/Vx1 current_steering_dac_unit_cell_with_encoder_19/Vbn
+ current_steering_dac_unit_cell_with_encoder_19/Vcn dummy_current_steering_dac_unit_cell_with_encoder_9/Vx1
+ current_steering_dac_unit_cell_with_encoder_6/I2 dummy_current_steering_dac_unit_cell_with_encoder_0/Vy
+ current_steering_dac_unit_cell_with_encoder_19/Vx current_steering_dac_unit_cell_with_encoder_6/I1
+ current_steering_dac_unit_cell_with_encoder_6/Vy current_steering_dac_unit_cell_with_encoder_19/VN2
+ current_steering_dac_unit_cell_with_encoder_9/Vbn current_steering_dac_unit_cell_with_encoder_9/Vcn
+ current_steering_dac_unit_cell_with_encoder_6/VP current_steering_dac_unit_cell_with_encoder_19/VP
+ dummy_current_steering_dac_unit_cell_with_encoder_9/VP dummy_current_steering_dac_unit_cell_with_encoder_3/Vx1
+ current_steering_dac_unit_cell_with_encoder_9/VN2 current_steering_dac_unit_cell_with_encoder_8/VP
+ current_steering_dac_unit_cell_with_encoder_8/Vx dummy_current_steering_dac_unit_cell_with_encoder_9/Vbn
+ dummy_current_steering_dac_unit_cell_with_encoder_9/I2 dummy_current_steering_dac_unit_cell_with_encoder_9/Vcn
+ current_steering_dac_unit_cell_with_encoder_8/I2 dummy_current_steering_dac_unit_cell_with_encoder_9/I1
+ current_steering_dac_unit_cell_with_encoder_8/I1 current_steering_dac_unit_cell_with_encoder_19/I2
+ dummy_current_steering_dac_unit_cell_with_encoder_9/Vy current_steering_dac_unit_cell_with_encoder_2/Vy
+ current_steering_dac_unit_cell_with_encoder_9/I2 dummy_current_steering_dac_unit_cell_with_encoder_9/VN2
+ current_steering_dac_unit_cell_with_encoder_19/I1 current_steering_dac_unit_cell_with_encoder_9/Vx
+ current_steering_dac_unit_cell_with_encoder_16/Vy current_steering_dac_unit_cell_with_encoder_9/I1
+ current_steering_dac_unit_cell_with_encoder_6/Vcn current_steering_dac_unit_cell_with_encoder_9/Vy
+ VSUBS current_steering_dac_unit_cell_with_encoder_6/Vx current_steering_dac_unit_cell_with_encoder_6/Vbn
Xdummy_current_steering_dac_unit_cell_with_encoder_0 current_steering_dac_unit_cell_with_encoder_19/I1
+ current_steering_dac_unit_cell_with_encoder_19/I2 current_steering_dac_unit_cell_with_encoder_19/Vbn
+ current_steering_dac_unit_cell_with_encoder_19/Vcn current_steering_dac_unit_cell_with_encoder_19/Vx
+ current_steering_dac_unit_cell_with_encoder_8/Vx dummy_current_steering_dac_unit_cell_with_encoder_0/Vy
+ current_steering_dac_unit_cell_with_encoder_19/VP VSUBS current_steering_dac_unit_cell_with_encoder_19/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_1 dummy_current_steering_dac_unit_cell_with_encoder_9/I1
+ dummy_current_steering_dac_unit_cell_with_encoder_9/I2 dummy_current_steering_dac_unit_cell_with_encoder_9/Vbn
+ dummy_current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx1
+ dummy_current_steering_dac_unit_cell_with_encoder_1/Vx1 current_steering_dac_unit_cell_with_encoder_16/Vy
+ dummy_current_steering_dac_unit_cell_with_encoder_9/VP VSUBS dummy_current_steering_dac_unit_cell_with_encoder_9/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_2 dummy_current_steering_dac_unit_cell_with_encoder_9/I1
+ dummy_current_steering_dac_unit_cell_with_encoder_9/I2 dummy_current_steering_dac_unit_cell_with_encoder_9/Vbn
+ dummy_current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx1
+ dummy_current_steering_dac_unit_cell_with_encoder_2/Vx1 current_steering_dac_unit_cell_with_encoder_9/Vy
+ dummy_current_steering_dac_unit_cell_with_encoder_9/VP VSUBS dummy_current_steering_dac_unit_cell_with_encoder_9/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_3 dummy_current_steering_dac_unit_cell_with_encoder_9/I1
+ dummy_current_steering_dac_unit_cell_with_encoder_9/I2 dummy_current_steering_dac_unit_cell_with_encoder_9/Vbn
+ dummy_current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx1
+ dummy_current_steering_dac_unit_cell_with_encoder_3/Vx1 current_steering_dac_unit_cell_with_encoder_6/Vy
+ dummy_current_steering_dac_unit_cell_with_encoder_9/VP VSUBS dummy_current_steering_dac_unit_cell_with_encoder_9/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_4 dummy_current_steering_dac_unit_cell_with_encoder_9/I1
+ dummy_current_steering_dac_unit_cell_with_encoder_9/I2 dummy_current_steering_dac_unit_cell_with_encoder_9/Vbn
+ dummy_current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx1
+ dummy_current_steering_dac_unit_cell_with_encoder_4/Vx1 current_steering_dac_unit_cell_with_encoder_2/Vy
+ dummy_current_steering_dac_unit_cell_with_encoder_9/VP VSUBS dummy_current_steering_dac_unit_cell_with_encoder_9/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_0 current_steering_dac_unit_cell_with_encoder_8/I1
+ current_steering_dac_unit_cell_with_encoder_8/I2 current_steering_dac_unit_cell_with_encoder_8/Vbn
+ current_steering_dac_unit_cell_with_encoder_8/Vcn current_steering_dac_unit_cell_with_encoder_8/Vx
+ current_steering_dac_unit_cell_with_encoder_9/Vx current_steering_dac_unit_cell_with_encoder_2/Vy
+ current_steering_dac_unit_cell_with_encoder_8/VP VSUBS current_steering_dac_unit_cell_with_encoder_8/VN2
+ current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_1 current_steering_dac_unit_cell_with_encoder_9/I1
+ current_steering_dac_unit_cell_with_encoder_9/I2 current_steering_dac_unit_cell_with_encoder_9/Vbn
+ current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_9/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx current_steering_dac_unit_cell_with_encoder_2/Vy
+ current_steering_dac_unit_cell_with_encoder_9/VP VSUBS current_steering_dac_unit_cell_with_encoder_9/VN2
+ current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_5 current_steering_dac_unit_cell_with_encoder_19/I1
+ current_steering_dac_unit_cell_with_encoder_19/I2 current_steering_dac_unit_cell_with_encoder_19/Vbn
+ current_steering_dac_unit_cell_with_encoder_19/Vcn current_steering_dac_unit_cell_with_encoder_19/Vx
+ current_steering_dac_unit_cell_with_encoder_8/Vx dummy_current_steering_dac_unit_cell_with_encoder_9/Vy
+ current_steering_dac_unit_cell_with_encoder_19/VP VSUBS current_steering_dac_unit_cell_with_encoder_19/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_2 current_steering_dac_unit_cell_with_encoder_6/I1
+ current_steering_dac_unit_cell_with_encoder_6/I2 current_steering_dac_unit_cell_with_encoder_6/Vbn
+ current_steering_dac_unit_cell_with_encoder_6/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx1 current_steering_dac_unit_cell_with_encoder_2/Vy
+ current_steering_dac_unit_cell_with_encoder_6/VP VSUBS current_steering_dac_unit_cell_with_encoder_6/VN2
+ current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_6 current_steering_dac_unit_cell_with_encoder_8/I1
+ current_steering_dac_unit_cell_with_encoder_8/I2 current_steering_dac_unit_cell_with_encoder_8/Vbn
+ current_steering_dac_unit_cell_with_encoder_8/Vcn current_steering_dac_unit_cell_with_encoder_8/Vx
+ current_steering_dac_unit_cell_with_encoder_9/Vx dummy_current_steering_dac_unit_cell_with_encoder_9/Vy
+ current_steering_dac_unit_cell_with_encoder_8/VP VSUBS current_steering_dac_unit_cell_with_encoder_8/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_7 current_steering_dac_unit_cell_with_encoder_9/I1
+ current_steering_dac_unit_cell_with_encoder_9/I2 current_steering_dac_unit_cell_with_encoder_9/Vbn
+ current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_9/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx dummy_current_steering_dac_unit_cell_with_encoder_9/Vy
+ current_steering_dac_unit_cell_with_encoder_9/VP VSUBS current_steering_dac_unit_cell_with_encoder_9/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_10 current_steering_dac_unit_cell_with_encoder_6/I1
+ current_steering_dac_unit_cell_with_encoder_6/I2 current_steering_dac_unit_cell_with_encoder_6/Vbn
+ current_steering_dac_unit_cell_with_encoder_6/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx1 current_steering_dac_unit_cell_with_encoder_9/Vy
+ current_steering_dac_unit_cell_with_encoder_6/VP VSUBS current_steering_dac_unit_cell_with_encoder_6/VN2
+ current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_4 current_steering_dac_unit_cell_with_encoder_8/I1
+ current_steering_dac_unit_cell_with_encoder_8/I2 current_steering_dac_unit_cell_with_encoder_8/Vbn
+ current_steering_dac_unit_cell_with_encoder_8/Vcn current_steering_dac_unit_cell_with_encoder_8/Vx
+ current_steering_dac_unit_cell_with_encoder_9/Vx current_steering_dac_unit_cell_with_encoder_6/Vy
+ current_steering_dac_unit_cell_with_encoder_8/VP VSUBS current_steering_dac_unit_cell_with_encoder_8/VN2
+ current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_8 current_steering_dac_unit_cell_with_encoder_6/I1
+ current_steering_dac_unit_cell_with_encoder_6/I2 current_steering_dac_unit_cell_with_encoder_6/Vbn
+ current_steering_dac_unit_cell_with_encoder_6/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx1 dummy_current_steering_dac_unit_cell_with_encoder_9/Vy
+ current_steering_dac_unit_cell_with_encoder_6/VP VSUBS current_steering_dac_unit_cell_with_encoder_6/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_5 current_steering_dac_unit_cell_with_encoder_9/I1
+ current_steering_dac_unit_cell_with_encoder_9/I2 current_steering_dac_unit_cell_with_encoder_9/Vbn
+ current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_9/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx current_steering_dac_unit_cell_with_encoder_6/Vy
+ current_steering_dac_unit_cell_with_encoder_9/VP VSUBS current_steering_dac_unit_cell_with_encoder_9/VN2
+ current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_9 dummy_current_steering_dac_unit_cell_with_encoder_9/I1
+ dummy_current_steering_dac_unit_cell_with_encoder_9/I2 dummy_current_steering_dac_unit_cell_with_encoder_9/Vbn
+ dummy_current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx1
+ dummy_current_steering_dac_unit_cell_with_encoder_9/Vx1 dummy_current_steering_dac_unit_cell_with_encoder_9/Vy
+ dummy_current_steering_dac_unit_cell_with_encoder_9/VP VSUBS dummy_current_steering_dac_unit_cell_with_encoder_9/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_13 current_steering_dac_unit_cell_with_encoder_9/I1
+ current_steering_dac_unit_cell_with_encoder_9/I2 current_steering_dac_unit_cell_with_encoder_9/Vbn
+ current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_9/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx current_steering_dac_unit_cell_with_encoder_16/Vy
+ current_steering_dac_unit_cell_with_encoder_9/VP VSUBS current_steering_dac_unit_cell_with_encoder_9/VN2
+ current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_12 current_steering_dac_unit_cell_with_encoder_8/I1
+ current_steering_dac_unit_cell_with_encoder_8/I2 current_steering_dac_unit_cell_with_encoder_8/Vbn
+ current_steering_dac_unit_cell_with_encoder_8/Vcn current_steering_dac_unit_cell_with_encoder_8/Vx
+ current_steering_dac_unit_cell_with_encoder_9/Vx current_steering_dac_unit_cell_with_encoder_16/Vy
+ current_steering_dac_unit_cell_with_encoder_8/VP VSUBS current_steering_dac_unit_cell_with_encoder_8/VN2
+ current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_6 current_steering_dac_unit_cell_with_encoder_6/I1
+ current_steering_dac_unit_cell_with_encoder_6/I2 current_steering_dac_unit_cell_with_encoder_6/Vbn
+ current_steering_dac_unit_cell_with_encoder_6/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx1 current_steering_dac_unit_cell_with_encoder_6/Vy
+ current_steering_dac_unit_cell_with_encoder_6/VP VSUBS current_steering_dac_unit_cell_with_encoder_6/VN2
+ current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_14 current_steering_dac_unit_cell_with_encoder_6/I1
+ current_steering_dac_unit_cell_with_encoder_6/I2 current_steering_dac_unit_cell_with_encoder_6/Vbn
+ current_steering_dac_unit_cell_with_encoder_6/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx1 current_steering_dac_unit_cell_with_encoder_16/Vy
+ current_steering_dac_unit_cell_with_encoder_6/VP VSUBS current_steering_dac_unit_cell_with_encoder_6/VN2
+ current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_9 current_steering_dac_unit_cell_with_encoder_9/I1
+ current_steering_dac_unit_cell_with_encoder_9/I2 current_steering_dac_unit_cell_with_encoder_9/Vbn
+ current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_9/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx current_steering_dac_unit_cell_with_encoder_9/Vy
+ current_steering_dac_unit_cell_with_encoder_9/VP VSUBS current_steering_dac_unit_cell_with_encoder_9/VN2
+ current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_8 current_steering_dac_unit_cell_with_encoder_8/I1
+ current_steering_dac_unit_cell_with_encoder_8/I2 current_steering_dac_unit_cell_with_encoder_8/Vbn
+ current_steering_dac_unit_cell_with_encoder_8/Vcn current_steering_dac_unit_cell_with_encoder_8/Vx
+ current_steering_dac_unit_cell_with_encoder_9/Vx current_steering_dac_unit_cell_with_encoder_9/Vy
+ current_steering_dac_unit_cell_with_encoder_8/VP VSUBS current_steering_dac_unit_cell_with_encoder_8/VN2
+ current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_16 current_steering_dac_unit_cell_with_encoder_19/I1
+ current_steering_dac_unit_cell_with_encoder_19/I2 current_steering_dac_unit_cell_with_encoder_19/Vbn
+ current_steering_dac_unit_cell_with_encoder_19/Vcn current_steering_dac_unit_cell_with_encoder_19/Vx
+ current_steering_dac_unit_cell_with_encoder_8/Vx current_steering_dac_unit_cell_with_encoder_16/Vy
+ current_steering_dac_unit_cell_with_encoder_19/VP VSUBS current_steering_dac_unit_cell_with_encoder_19/VN2
+ current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_10 current_steering_dac_unit_cell_with_encoder_8/I1
+ current_steering_dac_unit_cell_with_encoder_8/I2 current_steering_dac_unit_cell_with_encoder_8/Vbn
+ current_steering_dac_unit_cell_with_encoder_8/Vcn current_steering_dac_unit_cell_with_encoder_8/Vx
+ current_steering_dac_unit_cell_with_encoder_9/Vx dummy_current_steering_dac_unit_cell_with_encoder_0/Vy
+ current_steering_dac_unit_cell_with_encoder_8/VP VSUBS current_steering_dac_unit_cell_with_encoder_8/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_17 current_steering_dac_unit_cell_with_encoder_19/I1
+ current_steering_dac_unit_cell_with_encoder_19/I2 current_steering_dac_unit_cell_with_encoder_19/Vbn
+ current_steering_dac_unit_cell_with_encoder_19/Vcn current_steering_dac_unit_cell_with_encoder_19/Vx
+ current_steering_dac_unit_cell_with_encoder_8/Vx current_steering_dac_unit_cell_with_encoder_9/Vy
+ current_steering_dac_unit_cell_with_encoder_19/VP VSUBS current_steering_dac_unit_cell_with_encoder_19/VN2
+ current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_11 current_steering_dac_unit_cell_with_encoder_9/I1
+ current_steering_dac_unit_cell_with_encoder_9/I2 current_steering_dac_unit_cell_with_encoder_9/Vbn
+ current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_9/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx dummy_current_steering_dac_unit_cell_with_encoder_0/Vy
+ current_steering_dac_unit_cell_with_encoder_9/VP VSUBS current_steering_dac_unit_cell_with_encoder_9/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_18 current_steering_dac_unit_cell_with_encoder_19/I1
+ current_steering_dac_unit_cell_with_encoder_19/I2 current_steering_dac_unit_cell_with_encoder_19/Vbn
+ current_steering_dac_unit_cell_with_encoder_19/Vcn current_steering_dac_unit_cell_with_encoder_19/Vx
+ current_steering_dac_unit_cell_with_encoder_8/Vx current_steering_dac_unit_cell_with_encoder_6/Vy
+ current_steering_dac_unit_cell_with_encoder_19/VP VSUBS current_steering_dac_unit_cell_with_encoder_19/VN2
+ current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_12 current_steering_dac_unit_cell_with_encoder_6/I1
+ current_steering_dac_unit_cell_with_encoder_6/I2 current_steering_dac_unit_cell_with_encoder_6/Vbn
+ current_steering_dac_unit_cell_with_encoder_6/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx
+ current_steering_dac_unit_cell_with_encoder_6/Vx1 dummy_current_steering_dac_unit_cell_with_encoder_0/Vy
+ current_steering_dac_unit_cell_with_encoder_6/VP VSUBS current_steering_dac_unit_cell_with_encoder_6/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
Xcurrent_steering_dac_unit_cell_with_encoder_19 current_steering_dac_unit_cell_with_encoder_19/I1
+ current_steering_dac_unit_cell_with_encoder_19/I2 current_steering_dac_unit_cell_with_encoder_19/Vbn
+ current_steering_dac_unit_cell_with_encoder_19/Vcn current_steering_dac_unit_cell_with_encoder_19/Vx
+ current_steering_dac_unit_cell_with_encoder_8/Vx current_steering_dac_unit_cell_with_encoder_2/Vy
+ current_steering_dac_unit_cell_with_encoder_19/VP VSUBS current_steering_dac_unit_cell_with_encoder_19/VN2
+ current_steering_dac_unit_cell_with_encoder
Xdummy_current_steering_dac_unit_cell_with_encoder_13 dummy_current_steering_dac_unit_cell_with_encoder_9/I1
+ dummy_current_steering_dac_unit_cell_with_encoder_9/I2 dummy_current_steering_dac_unit_cell_with_encoder_9/Vbn
+ dummy_current_steering_dac_unit_cell_with_encoder_9/Vcn current_steering_dac_unit_cell_with_encoder_6/Vx1
+ dummy_current_steering_dac_unit_cell_with_encoder_13/Vx1 dummy_current_steering_dac_unit_cell_with_encoder_0/Vy
+ dummy_current_steering_dac_unit_cell_with_encoder_9/VP VSUBS dummy_current_steering_dac_unit_cell_with_encoder_9/VN2
+ dummy_current_steering_dac_unit_cell_with_encoder
.ends

**.subckt current_steering_dac X0 X1 X2 X3 Y0 Y1 Y2 Y3 I1 I2 VDD GND Vbn Vcn
Xhalf_dac_for_mirroring_1 GND GND GND GND Vbn Vcn GND VDD GND GND Vbn Vcn GND I2 GND
+ X0 I1 Y1 GND Vbn Vcn VDD VDD VDD GND GND VDD X1 Vbn I2 Vcn I2 I1 I1 I2 GND Y0 I2
+ GND I1 X2 Y3 I1 Vcn Y2 GND X3 Vbn half_dac_for_mirroring
Xhalf_dac_for_mirroring_0 GND GND GND GND Vbn Vcn GND VDD GND GND Vbn Vcn GND I2 GND
+ X0 I1 Y1 GND Vbn Vcn VDD VDD VDD GND GND VDD X1 Vbn I2 Vcn I2 I1 I1 I2 GND Y0 I2
+ GND I1 X2 Y3 I1 Vcn Y2 GND X3 Vbn half_dac_for_mirroring
**.ends

