magic
tech sky130A
timestamp 1702417875
<< locali >>
rect -2520 8215 -2480 8225
rect -2520 8195 -2510 8215
rect -2490 8195 -2480 8215
rect -2520 8100 -2480 8195
rect -1870 8215 -1830 8225
rect -1870 8195 -1860 8215
rect -1840 8195 -1830 8215
rect -2520 8080 -2510 8100
rect -2490 8080 -2480 8100
rect -2520 8070 -2480 8080
rect -2090 7970 -2070 8110
rect -2050 8030 -2030 8110
rect -2010 8070 -1990 8110
rect -1970 8090 -1930 8110
rect -2010 8050 -1970 8070
rect -2050 8020 -2010 8030
rect -2050 8000 -2040 8020
rect -2020 8000 -2010 8020
rect -2050 7990 -2010 8000
rect -1990 8010 -1970 8050
rect -1950 8050 -1930 8090
rect -1870 8100 -1830 8195
rect -1220 8215 -1180 8225
rect -1220 8195 -1210 8215
rect -1190 8195 -1180 8215
rect -1870 8080 -1860 8100
rect -1840 8080 -1830 8100
rect -1870 8070 -1830 8080
rect -1560 8090 -1320 8110
rect -1560 8050 -1540 8090
rect -1400 8060 -1360 8070
rect -1400 8050 -1390 8060
rect -1950 8030 -1540 8050
rect -1520 8040 -1390 8050
rect -1370 8040 -1360 8060
rect -1520 8030 -1360 8040
rect -1340 8050 -1320 8090
rect -1220 8100 -1180 8195
rect -570 8215 -530 8225
rect -570 8195 -560 8215
rect -540 8195 -530 8215
rect -1220 8080 -1210 8100
rect -1190 8080 -1180 8100
rect -1220 8070 -1180 8080
rect -910 8100 -710 8110
rect -910 8090 -740 8100
rect -910 8050 -890 8090
rect -750 8080 -740 8090
rect -720 8080 -710 8100
rect -750 8070 -710 8080
rect -570 8100 -530 8195
rect -570 8080 -560 8100
rect -540 8080 -530 8100
rect -570 8070 -530 8080
rect 1030 8215 1070 8225
rect 1030 8195 1040 8215
rect 1060 8195 1070 8215
rect 1030 8100 1070 8195
rect 1030 8080 1040 8100
rect 1060 8080 1070 8100
rect 1030 8070 1070 8080
rect 1680 8215 1720 8225
rect 1680 8195 1690 8215
rect 1710 8195 1720 8215
rect 1680 8100 1720 8195
rect 1680 8080 1690 8100
rect 1710 8080 1720 8100
rect 1680 8070 1720 8080
rect 2330 8215 2370 8225
rect 2330 8195 2340 8215
rect 2360 8195 2370 8215
rect 2330 8100 2370 8195
rect 2330 8080 2340 8100
rect 2360 8080 2370 8100
rect 2330 8070 2370 8080
rect 2980 8215 3020 8225
rect 2980 8195 2990 8215
rect 3010 8195 3020 8215
rect 2980 8100 3020 8195
rect 2980 8080 2990 8100
rect 3010 8080 3020 8100
rect 2980 8070 3020 8080
rect -1340 8030 -890 8050
rect -870 8030 140 8050
rect -1520 8010 -1500 8030
rect -870 8010 -850 8030
rect 120 8010 140 8030
rect -1990 7990 -1500 8010
rect -1480 7990 -850 8010
rect -830 7990 100 8010
rect 120 7990 710 8010
rect -1480 7970 -1460 7990
rect -830 7970 -810 7990
rect 80 7970 100 7990
rect 690 7970 710 7990
rect -2090 7950 -1460 7970
rect -1440 7950 -810 7970
rect -790 7950 60 7970
rect 80 7950 670 7970
rect 690 7950 1320 7970
rect -2090 7930 -2070 7950
rect -1440 7930 -1420 7950
rect -790 7930 -770 7950
rect 40 7930 60 7950
rect 650 7930 670 7950
rect 1300 7930 1320 7950
rect -3350 7920 -3310 7930
rect -3350 7900 -3340 7920
rect -3320 7900 -3310 7920
rect -3350 7890 -3310 7900
rect -2700 7920 -2070 7930
rect -2700 7900 -2690 7920
rect -2670 7910 -2070 7920
rect -2050 7920 -1420 7930
rect -2670 7900 -2660 7910
rect -2700 7890 -2660 7900
rect -2050 7900 -2040 7920
rect -2020 7910 -1420 7920
rect -1400 7920 -770 7930
rect -2020 7900 -2010 7910
rect -2050 7890 -2010 7900
rect -1400 7900 -1390 7920
rect -1370 7910 -770 7920
rect -750 7920 20 7930
rect -1370 7900 -1360 7910
rect -1400 7890 -1360 7900
rect -750 7900 -740 7920
rect -720 7910 20 7920
rect 40 7910 630 7930
rect 650 7910 1280 7930
rect 1300 7910 1930 7930
rect -720 7900 -710 7910
rect -750 7890 -710 7900
rect 0 7890 20 7910
rect 610 7890 630 7910
rect 1260 7890 1280 7910
rect 1910 7890 1930 7910
rect -130 7810 0 7830
rect -130 6655 -110 7810
rect -150 6635 -110 6655
rect -40 6520 0 6530
rect -40 6500 -30 6520
rect -10 6500 0 6520
rect -40 6490 0 6500
rect -150 5330 -95 5340
rect -150 5320 -125 5330
rect -135 5310 -125 5320
rect -105 5310 -95 5330
rect -135 5300 -95 5310
rect -135 5190 0 5200
rect -135 5170 -125 5190
rect -105 5180 0 5190
rect -105 5170 -95 5180
rect -135 5160 -95 5170
rect -150 4005 -110 4025
rect -130 3885 -110 4005
rect -130 3865 0 3885
rect -135 2720 -95 2730
rect -135 2710 -125 2720
rect -150 2700 -125 2710
rect -105 2700 -95 2720
rect -150 2690 -95 2700
rect -95 2580 -55 2590
rect -95 2560 -85 2580
rect -65 2570 -55 2580
rect -65 2560 0 2570
rect -95 2550 0 2560
rect -65 1405 -25 1415
rect -65 1395 -55 1405
rect -150 1385 -55 1395
rect -35 1385 -25 1405
rect -150 1375 -25 1385
rect -130 1235 0 1255
rect -130 80 -110 1235
rect -150 60 -110 80
<< viali >>
rect -2510 8195 -2490 8215
rect -1860 8195 -1840 8215
rect -2510 8080 -2490 8100
rect -2040 8000 -2020 8020
rect -1210 8195 -1190 8215
rect -1860 8080 -1840 8100
rect -1390 8040 -1370 8060
rect -560 8195 -540 8215
rect -1210 8080 -1190 8100
rect -740 8080 -720 8100
rect -560 8080 -540 8100
rect 1040 8195 1060 8215
rect 1040 8080 1060 8100
rect 1690 8195 1710 8215
rect 1690 8080 1710 8100
rect 2340 8195 2360 8215
rect 2340 8080 2360 8100
rect 2990 8195 3010 8215
rect 2990 8080 3010 8100
rect -3340 7900 -3320 7920
rect -2690 7900 -2670 7920
rect -2040 7900 -2020 7920
rect -1390 7900 -1370 7920
rect -740 7900 -720 7920
rect -30 6500 -10 6520
rect -125 5310 -105 5330
rect -125 5170 -105 5190
rect -125 2700 -105 2720
rect -85 2560 -65 2580
rect -55 1385 -35 1405
<< metal1 >>
rect -2520 8215 -2480 8225
rect -1870 8215 -1830 8225
rect -1220 8215 -1180 8225
rect -570 8215 -530 8225
rect 1030 8215 1070 8225
rect 1680 8215 1720 8225
rect 2330 8215 2370 8225
rect 2980 8215 3020 8225
rect -3165 8195 -2510 8215
rect -2490 8195 -1860 8215
rect -1840 8195 -1210 8215
rect -1190 8195 -560 8215
rect -540 8195 1040 8215
rect 1060 8195 1690 8215
rect 1710 8195 2340 8215
rect 2360 8195 2990 8215
rect 3010 8195 3365 8215
rect -3165 8185 3365 8195
rect -3350 7920 -3310 7930
rect -3350 7900 -3340 7920
rect -3320 7900 -3310 7920
rect -3350 7890 -3310 7900
rect -3165 7890 -3135 8185
rect -2950 8125 3365 8155
rect -2950 7890 -2920 8125
rect -2520 8100 -2480 8110
rect -2520 8080 -2510 8100
rect -2490 8080 -2480 8100
rect -2520 8070 -2480 8080
rect -2700 7920 -2660 7930
rect -2700 7900 -2690 7920
rect -2670 7900 -2660 7920
rect -2700 7890 -2660 7900
rect -2515 7890 -2485 8070
rect -2300 7890 -2270 8125
rect -1870 8100 -1830 8110
rect -1870 8080 -1860 8100
rect -1840 8080 -1830 8100
rect -1870 8070 -1830 8080
rect -2050 8020 -2010 8030
rect -2050 8000 -2040 8020
rect -2020 8000 -2010 8020
rect -2050 7990 -2010 8000
rect -2025 7930 -2010 7990
rect -2050 7920 -2010 7930
rect -2050 7900 -2040 7920
rect -2020 7900 -2010 7920
rect -2050 7890 -2010 7900
rect -1865 7890 -1835 8070
rect -1650 7890 -1620 8125
rect -1220 8100 -1180 8110
rect -1220 8080 -1210 8100
rect -1190 8080 -1180 8100
rect -1220 8070 -1180 8080
rect -1400 8060 -1360 8070
rect -1400 8040 -1390 8060
rect -1370 8040 -1360 8060
rect -1400 8030 -1360 8040
rect -1375 7930 -1360 8030
rect -1400 7920 -1360 7930
rect -1400 7900 -1390 7920
rect -1370 7900 -1360 7920
rect -1400 7890 -1360 7900
rect -1215 7890 -1185 8070
rect -1000 7890 -970 8125
rect -750 8100 -710 8110
rect -750 8080 -740 8100
rect -720 8080 -710 8100
rect -750 8070 -710 8080
rect -570 8100 -530 8110
rect -570 8080 -560 8100
rect -540 8080 -530 8100
rect -570 8070 -530 8080
rect -725 7930 -710 8070
rect -750 7920 -710 7930
rect -750 7900 -740 7920
rect -720 7900 -710 7920
rect -750 7890 -710 7900
rect -565 7890 -535 8070
rect -350 7890 -320 8125
rect 170 7890 200 8125
rect 820 7890 850 8125
rect 1030 8100 1070 8110
rect 1030 8080 1040 8100
rect 1060 8080 1070 8100
rect 1030 8070 1070 8080
rect 1035 7890 1065 8070
rect 1470 7890 1500 8125
rect 1680 8100 1720 8110
rect 1680 8080 1690 8100
rect 1710 8080 1720 8100
rect 1680 8070 1720 8080
rect 1685 7890 1715 8070
rect 2120 7890 2150 8125
rect 2330 8100 2370 8110
rect 2330 8080 2340 8100
rect 2360 8080 2370 8100
rect 2330 8070 2370 8080
rect 2335 7890 2365 8070
rect 2770 7890 2800 8125
rect 2980 8100 3020 8110
rect 2980 8080 2990 8100
rect 3010 8080 3020 8100
rect 2980 8070 3020 8080
rect 2985 7890 3015 8070
rect -40 6520 0 6530
rect -40 6500 -30 6520
rect -10 6500 0 6520
rect -40 6490 0 6500
rect -135 5330 -95 5340
rect -135 5310 -125 5330
rect -105 5315 -95 5330
rect -105 5310 -65 5315
rect -135 5300 -65 5310
rect -135 5190 -95 5200
rect -135 5170 -125 5190
rect -105 5170 -95 5190
rect -135 5160 -95 5170
rect -135 2730 -120 5160
rect -135 2720 -95 2730
rect -135 2700 -125 2720
rect -105 2700 -95 2720
rect -135 2690 -95 2700
rect -80 2590 -65 5300
rect -95 2580 -55 2590
rect -95 2560 -85 2580
rect -65 2560 -55 2580
rect -95 2550 -55 2560
rect -40 1415 -25 6490
rect -65 1405 -25 1415
rect -65 1385 -55 1405
rect -35 1385 -25 1405
rect -65 1375 -25 1385
use half_dac_for_mirroring  half_dac_for_mirroring_0
timestamp 1702367632
transform 1 0 650 0 1 1315
box -650 -1315 2600 6575
use half_dac_for_mirroring  half_dac_for_mirroring_1
timestamp 1702367632
transform -1 0 -800 0 -1 6575
box -650 -1315 2600 6575
<< end >>
