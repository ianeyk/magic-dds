magic
tech sky130A
timestamp 1702595941
<< error_s >>
rect -236 5740 -235 5746
rect 414 5740 415 5746
rect 1064 5740 1065 5746
rect 1714 5740 1715 5746
rect 2364 5740 2365 5746
rect -230 5734 -224 5735
rect 420 5734 426 5735
rect 1070 5734 1076 5735
rect 1720 5734 1726 5735
rect 2370 5734 2376 5735
rect 2364 4425 2365 4431
rect 2370 4419 2376 4420
rect 2364 3110 2365 3116
rect 2370 3104 2376 3105
rect 2364 1795 2365 1801
rect 2370 1789 2376 1790
rect 2364 480 2365 486
rect 2370 474 2376 475
rect -236 -835 -235 -829
rect 414 -835 415 -829
rect 1064 -835 1065 -829
rect 1714 -835 1715 -829
rect 2364 -835 2365 -829
rect -230 -841 -224 -840
rect 420 -841 426 -840
rect 1070 -841 1076 -840
rect 1720 -841 1726 -840
rect 2370 -841 2376 -840
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_0
timestamp 1702593820
transform 1 0 0 0 1 15
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_1
timestamp 1702593820
transform 1 0 650 0 1 15
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_2
timestamp 1702593820
transform 1 0 1300 0 1 15
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_4
timestamp 1702593820
transform 1 0 0 0 1 1330
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_5
timestamp 1702593820
transform 1 0 650 0 1 1330
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_6
timestamp 1702593820
transform 1 0 1300 0 1 1330
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_8
timestamp 1702593820
transform 1 0 0 0 1 2645
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_9
timestamp 1702593820
transform 1 0 650 0 1 2645
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_10
timestamp 1702593820
transform 1 0 1300 0 1 2645
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_12
timestamp 1702593820
transform 1 0 0 0 1 3960
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_13
timestamp 1702593820
transform 1 0 650 0 1 3960
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_14
timestamp 1702593820
transform 1 0 1300 0 1 3960
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_16
timestamp 1702593820
transform 1 0 -650 0 1 3960
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_17
timestamp 1702593820
transform 1 0 -650 0 1 2645
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_18
timestamp 1702593820
transform 1 0 -650 0 1 1330
box 0 -15 650 1300
use current_steering_dac_unit_cell_with_encoder  current_steering_dac_unit_cell_with_encoder_19
timestamp 1702593820
transform 1 0 -650 0 1 15
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_0 ~/dev/git/magic-dds/magic
timestamp 1702591987
transform 1 0 -650 0 1 5275
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_1
timestamp 1702591987
transform 1 0 1950 0 1 3960
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_2
timestamp 1702591987
transform 1 0 1950 0 1 2645
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_3
timestamp 1702591987
transform 1 0 1950 0 1 1330
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_4
timestamp 1702591987
transform 1 0 1950 0 1 15
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_5
timestamp 1702591987
transform 1 0 -650 0 1 -1300
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_6
timestamp 1702591987
transform 1 0 0 0 1 -1300
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_7
timestamp 1702591987
transform 1 0 650 0 1 -1300
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_8
timestamp 1702591987
transform 1 0 1300 0 1 -1300
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_9
timestamp 1702591987
transform 1 0 1950 0 1 -1300
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_10
timestamp 1702591987
transform 1 0 0 0 1 5275
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_11
timestamp 1702591987
transform 1 0 650 0 1 5275
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_12
timestamp 1702591987
transform 1 0 1300 0 1 5275
box 0 -15 650 1300
use dummy_current_steering_dac_unit_cell_with_encoder  dummy_current_steering_dac_unit_cell_with_encoder_13
timestamp 1702591987
transform 1 0 1950 0 1 5275
box 0 -15 650 1300
<< end >>
