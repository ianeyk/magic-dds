magic
tech sky130A
timestamp 1702798187
<< nwell >>
rect -20 615 200 1675
<< nmos >>
rect 50 0 65 400
rect 115 0 130 400
<< pmos >>
rect 50 635 65 1655
rect 115 635 130 1655
<< ndiff >>
rect 0 385 50 400
rect 0 15 15 385
rect 35 15 50 385
rect 0 0 50 15
rect 65 385 115 400
rect 65 15 80 385
rect 100 15 115 385
rect 65 0 115 15
rect 130 385 180 400
rect 130 15 145 385
rect 165 15 180 385
rect 130 0 180 15
<< pdiff >>
rect 0 1640 50 1655
rect 0 645 15 1640
rect 35 645 50 1640
rect 0 635 50 645
rect 65 1640 115 1655
rect 65 645 80 1640
rect 100 645 115 1640
rect 65 635 115 645
rect 130 1640 180 1655
rect 130 645 145 1640
rect 165 645 180 1640
rect 130 635 180 645
<< ndiffc >>
rect 15 15 35 385
rect 80 15 100 385
rect 145 15 165 385
<< pdiffc >>
rect 15 645 35 1640
rect 80 645 100 1640
rect 145 645 165 1640
<< poly >>
rect 35 1700 75 1710
rect 35 1680 45 1700
rect 65 1680 75 1700
rect 35 1670 75 1680
rect 105 1700 145 1710
rect 105 1680 115 1700
rect 135 1680 145 1700
rect 105 1670 145 1680
rect 50 1655 65 1670
rect 115 1655 130 1670
rect 50 495 65 635
rect 115 560 130 635
rect 90 550 130 560
rect 90 530 100 550
rect 120 530 130 550
rect 90 520 130 530
rect 50 480 130 495
rect 50 445 90 455
rect 50 425 60 445
rect 80 425 90 445
rect 50 415 90 425
rect 50 400 65 415
rect 115 400 130 480
rect 50 -15 65 0
rect 115 -15 130 0
<< polycont >>
rect 45 1680 65 1700
rect 115 1680 135 1700
rect 100 530 120 550
rect 60 425 80 445
<< locali >>
rect 35 1700 75 1710
rect 35 1680 45 1700
rect 65 1680 75 1700
rect 35 1670 75 1680
rect 105 1700 145 1710
rect 105 1680 115 1700
rect 135 1680 145 1700
rect 105 1670 145 1680
rect 5 1640 45 1650
rect 5 645 15 1640
rect 35 645 45 1640
rect 5 475 45 645
rect 70 1640 110 1650
rect 70 645 80 1640
rect 100 645 110 1640
rect 70 610 110 645
rect 70 590 80 610
rect 100 590 110 610
rect 70 580 110 590
rect 135 1640 175 1650
rect 135 645 145 1640
rect 165 645 175 1640
rect 135 580 175 645
rect 70 550 130 560
rect 70 530 100 550
rect 120 530 130 550
rect 70 520 130 530
rect 5 395 30 475
rect 70 455 110 520
rect 150 500 175 580
rect 50 445 110 455
rect 50 425 60 445
rect 80 425 110 445
rect 50 415 110 425
rect 5 385 45 395
rect 5 15 15 385
rect 35 15 45 385
rect 5 5 45 15
rect 70 385 110 395
rect 70 15 80 385
rect 100 15 110 385
rect 70 5 110 15
rect 135 385 175 500
rect 135 15 145 385
rect 165 15 175 385
rect 135 5 175 15
<< viali >>
rect 80 590 100 610
rect 80 365 100 385
<< metal1 >>
rect 70 610 110 620
rect 70 590 80 610
rect 100 590 110 610
rect 70 385 110 590
rect 70 365 80 385
rect 100 365 110 385
rect 70 355 110 365
<< labels >>
flabel locali 55 1710 55 1710 1 FreeSans 160 0 0 0 phi1
port 1 n
flabel locali 125 1710 125 1710 1 FreeSans 160 0 0 0 phi2
port 2 n
<< end >>
