magic
tech sky130A
timestamp 1702624015
<< nwell >>
rect -130 130 800 270
<< nmos >>
rect 20 -5 35 95
rect 85 -5 100 95
rect 230 -5 245 95
rect 295 -5 310 95
rect 440 -5 455 95
rect 505 -5 520 95
rect 650 -5 665 95
rect 715 -5 730 95
<< pmos >>
rect 20 150 35 250
rect 85 150 100 250
rect 230 150 245 250
rect 295 150 310 250
rect 440 150 455 250
rect 505 150 520 250
rect 650 150 665 250
rect 715 150 730 250
<< ndiff >>
rect -30 80 20 95
rect -30 10 -15 80
rect 5 10 20 80
rect -30 -5 20 10
rect 35 80 85 95
rect 35 10 50 80
rect 70 10 85 80
rect 35 -5 85 10
rect 100 80 150 95
rect 100 10 115 80
rect 135 10 150 80
rect 100 -5 150 10
rect 180 80 230 95
rect 180 10 195 80
rect 215 10 230 80
rect 180 -5 230 10
rect 245 80 295 95
rect 245 10 260 80
rect 280 10 295 80
rect 245 -5 295 10
rect 310 80 360 95
rect 310 10 325 80
rect 345 10 360 80
rect 310 -5 360 10
rect 390 80 440 95
rect 390 10 405 80
rect 425 10 440 80
rect 390 -5 440 10
rect 455 80 505 95
rect 455 10 470 80
rect 490 10 505 80
rect 455 -5 505 10
rect 520 80 570 95
rect 520 10 535 80
rect 555 10 570 80
rect 520 -5 570 10
rect 600 80 650 95
rect 600 10 615 80
rect 635 10 650 80
rect 600 -5 650 10
rect 665 -5 715 95
rect 730 80 780 95
rect 730 10 745 80
rect 765 10 780 80
rect 730 -5 780 10
<< pdiff >>
rect -30 235 20 250
rect -30 165 -15 235
rect 5 165 20 235
rect -30 150 20 165
rect 35 150 85 250
rect 100 235 150 250
rect 100 165 115 235
rect 135 165 150 235
rect 100 150 150 165
rect 180 235 230 250
rect 180 165 195 235
rect 215 165 230 235
rect 180 150 230 165
rect 245 235 295 250
rect 245 165 260 235
rect 280 165 295 235
rect 245 150 295 165
rect 310 235 360 250
rect 310 165 325 235
rect 345 165 360 235
rect 310 150 360 165
rect 390 235 440 250
rect 390 165 405 235
rect 425 165 440 235
rect 390 150 440 165
rect 455 235 505 250
rect 455 165 470 235
rect 490 165 505 235
rect 455 150 505 165
rect 520 235 570 250
rect 520 165 535 235
rect 555 165 570 235
rect 520 150 570 165
rect 600 235 650 250
rect 600 165 615 235
rect 635 165 650 235
rect 600 150 650 165
rect 665 235 715 250
rect 665 165 680 235
rect 700 165 715 235
rect 665 150 715 165
rect 730 235 780 250
rect 730 165 745 235
rect 765 165 780 235
rect 730 150 780 165
<< ndiffc >>
rect -15 10 5 80
rect 50 10 70 80
rect 115 10 135 80
rect 195 10 215 80
rect 260 10 280 80
rect 325 10 345 80
rect 405 10 425 80
rect 470 10 490 80
rect 535 10 555 80
rect 615 10 635 80
rect 745 10 765 80
<< pdiffc >>
rect -15 165 5 235
rect 115 165 135 235
rect 195 165 215 235
rect 260 165 280 235
rect 325 165 345 235
rect 405 165 425 235
rect 470 165 490 235
rect 535 165 555 235
rect 615 165 635 235
rect 680 165 700 235
rect 745 165 765 235
<< psubdiff >>
rect -110 80 -60 95
rect -110 10 -95 80
rect -75 10 -60 80
rect -110 -5 -60 10
<< nsubdiff >>
rect -110 235 -60 250
rect -110 165 -95 235
rect -75 165 -60 235
rect -110 150 -60 165
<< psubdiffcont >>
rect -95 10 -75 80
<< nsubdiffcont >>
rect -95 165 -75 235
<< poly >>
rect 285 435 325 445
rect 285 415 295 435
rect 315 415 325 435
rect 285 405 325 415
rect 295 345 310 405
rect -5 335 35 345
rect -5 315 5 335
rect 25 315 35 335
rect -5 305 35 315
rect 20 250 35 305
rect 85 335 125 345
rect 85 315 95 335
rect 115 315 125 335
rect 85 305 125 315
rect 285 335 325 345
rect 285 315 295 335
rect 315 315 325 335
rect 285 305 325 315
rect 625 335 665 345
rect 625 315 635 335
rect 655 315 665 335
rect 625 305 665 315
rect 85 250 100 305
rect 205 295 245 305
rect 205 275 215 295
rect 235 275 245 295
rect 205 265 245 275
rect 230 250 245 265
rect 295 250 310 305
rect 415 295 455 305
rect 415 275 425 295
rect 445 275 455 295
rect 415 265 455 275
rect 440 250 455 265
rect 505 295 545 305
rect 505 275 515 295
rect 535 275 545 295
rect 505 265 545 275
rect 505 250 520 265
rect 650 250 665 305
rect 715 335 755 345
rect 715 315 725 335
rect 745 315 755 335
rect 715 305 755 315
rect 715 250 730 305
rect 20 95 35 150
rect 85 95 100 150
rect 230 95 245 150
rect 295 95 310 150
rect 440 95 455 150
rect 505 95 520 150
rect 650 95 665 150
rect 715 95 730 150
rect 20 -20 35 -5
rect 85 -20 100 -5
rect 230 -20 245 -5
rect 295 -20 310 -5
rect 440 -20 455 -5
rect 505 -20 520 -5
rect 650 -20 665 -5
rect 715 -20 730 -5
<< polycont >>
rect 295 415 315 435
rect 5 315 25 335
rect 95 315 115 335
rect 295 315 315 335
rect 635 315 655 335
rect 215 275 235 295
rect 425 275 445 295
rect 515 275 535 295
rect 725 315 745 335
<< locali >>
rect 15 385 35 445
rect 285 435 325 445
rect 285 415 295 435
rect 315 415 325 435
rect 285 405 325 415
rect 15 365 735 385
rect 15 345 35 365
rect 715 345 735 365
rect -5 335 35 345
rect -5 315 5 335
rect 25 315 35 335
rect -5 305 35 315
rect 85 335 665 345
rect 85 315 95 335
rect 115 325 295 335
rect 115 315 125 325
rect 85 305 125 315
rect 285 315 295 325
rect 315 325 635 335
rect 315 315 325 325
rect 285 305 325 315
rect 625 315 635 325
rect 655 315 665 335
rect 625 305 665 315
rect 715 335 755 345
rect 715 315 725 335
rect 745 315 755 335
rect 715 305 755 315
rect 205 295 245 305
rect 205 285 215 295
rect -5 275 215 285
rect 235 275 245 295
rect 415 295 455 305
rect 415 285 425 295
rect -5 265 245 275
rect 335 275 425 285
rect 445 275 455 295
rect 335 265 455 275
rect 505 295 545 305
rect 505 275 515 295
rect 535 285 545 295
rect 535 275 755 285
rect 505 265 755 275
rect -5 245 15 265
rect 335 245 355 265
rect 605 245 625 265
rect 735 245 755 265
rect -105 235 -65 245
rect -105 175 -95 235
rect -145 165 -95 175
rect -75 165 -65 235
rect -145 155 -65 165
rect -25 235 15 245
rect -25 165 -15 235
rect 5 165 15 235
rect -25 155 15 165
rect 105 235 145 245
rect 105 165 115 235
rect 135 165 145 235
rect 105 155 145 165
rect 185 235 225 245
rect 185 165 195 235
rect 215 165 225 235
rect 185 155 225 165
rect 250 235 290 245
rect 250 165 260 235
rect 280 165 290 235
rect 250 155 290 165
rect 315 235 355 245
rect 315 165 325 235
rect 345 165 355 235
rect 315 155 355 165
rect 395 235 435 245
rect 395 165 405 235
rect 425 165 435 235
rect 395 155 435 165
rect 460 235 500 245
rect 460 165 470 235
rect 490 165 500 235
rect 460 155 500 165
rect 525 235 565 245
rect 525 165 535 235
rect 555 165 565 235
rect 525 155 565 165
rect 605 235 645 245
rect 605 165 615 235
rect 635 165 645 235
rect 605 155 645 165
rect 670 235 710 245
rect 670 165 680 235
rect 700 165 710 235
rect 670 155 710 165
rect 735 235 775 245
rect 735 165 745 235
rect 765 165 775 235
rect 735 155 775 165
rect -145 -15 -125 155
rect -5 130 15 155
rect -5 110 125 130
rect -5 90 15 110
rect 105 90 125 110
rect 195 90 215 155
rect 325 90 345 155
rect 405 90 425 155
rect 535 90 555 155
rect 745 90 765 155
rect -105 80 -65 90
rect -105 10 -95 80
rect -75 10 -65 80
rect -105 0 -65 10
rect -25 80 15 90
rect -25 10 -15 80
rect 5 10 15 80
rect -25 0 15 10
rect 40 80 80 90
rect 40 10 50 80
rect 70 10 80 80
rect 40 0 80 10
rect 105 80 145 90
rect 105 10 115 80
rect 135 10 145 80
rect 105 0 145 10
rect 185 80 225 90
rect 185 10 195 80
rect 215 10 225 80
rect 185 0 225 10
rect 250 80 290 90
rect 250 10 260 80
rect 280 10 290 80
rect 250 0 290 10
rect 315 80 355 90
rect 315 10 325 80
rect 345 10 355 80
rect 315 0 355 10
rect 395 80 435 90
rect 395 10 405 80
rect 425 10 435 80
rect 395 0 435 10
rect 460 80 500 90
rect 460 10 470 80
rect 490 10 500 80
rect 460 0 500 10
rect 525 80 565 90
rect 525 10 535 80
rect 555 10 565 80
rect 525 0 565 10
rect 605 80 645 90
rect 605 10 615 80
rect 635 10 645 80
rect 605 0 645 10
rect 735 80 775 90
rect 735 10 745 80
rect 765 10 775 80
rect 735 0 775 10
rect 195 -20 215 0
rect 405 -20 425 0
rect 535 -20 555 0
<< viali >>
rect -95 165 -75 235
rect 115 165 135 235
rect 260 165 280 235
rect 470 165 490 235
rect 680 165 700 235
rect -95 10 -75 80
rect 50 10 70 80
rect 260 10 280 80
rect 470 10 490 80
rect 615 10 635 80
<< metal1 >>
rect -145 235 800 250
rect -145 165 -95 235
rect -75 165 115 235
rect 135 165 260 235
rect 280 165 470 235
rect 490 165 680 235
rect 700 165 800 235
rect -145 150 800 165
rect -145 80 800 95
rect -145 10 -95 80
rect -75 10 50 80
rect 70 10 260 80
rect 280 10 470 80
rect 490 10 615 80
rect 635 10 800 80
rect -145 -5 800 10
<< labels >>
flabel locali 25 445 25 445 1 FreeSans 160 0 0 0 b0
port 1 n
flabel locali 305 445 305 445 1 FreeSans 160 0 0 0 b1
port 2 n
flabel locali 205 -20 205 -20 5 FreeSans 160 0 0 0 y1
port 4 s
flabel locali 415 -20 415 -20 5 FreeSans 160 0 0 0 y2
port 5 s
flabel locali 545 -20 545 -20 5 FreeSans 160 0 0 0 y3
port 6 s
flabel metal1 -145 200 -145 200 7 FreeSans 160 0 0 0 VP
port 7 w
flabel metal1 -145 45 -145 45 7 FreeSans 160 0 0 0 VN
port 8 w
<< end >>
