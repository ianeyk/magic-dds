magic
tech sky130A
timestamp 1702617854
<< nwell >>
rect -70 375 1340 2160
<< nmos >>
rect 0 40 50 340
rect 100 40 150 340
rect 280 40 330 340
rect 380 40 430 340
rect 560 40 610 340
rect 660 40 710 340
rect 840 40 890 340
rect 940 40 990 340
rect 1120 40 1170 340
rect 1220 40 1270 340
rect 160 -370 210 -70
rect 260 -370 310 -70
rect 360 -370 410 -70
rect 460 -370 510 -70
rect 560 -370 610 -70
rect 660 -370 710 -70
rect 760 -370 810 -70
rect 860 -370 910 -70
rect 960 -370 1010 -70
rect 1060 -370 1110 -70
<< pmos >>
rect 160 1340 210 2140
rect 260 1340 310 2140
rect 360 1340 410 2140
rect 460 1340 510 2140
rect 560 1340 610 2140
rect 660 1340 710 2140
rect 760 1340 810 2140
rect 860 1340 910 2140
rect 960 1340 1010 2140
rect 1060 1340 1110 2140
rect 0 395 50 1195
rect 100 395 150 1195
rect 280 395 330 1195
rect 380 395 430 1195
rect 560 395 610 1195
rect 660 395 710 1195
rect 840 395 890 1195
rect 940 395 990 1195
rect 1120 395 1170 1195
rect 1220 395 1270 1195
<< ndiff >>
rect -50 325 0 340
rect -50 55 -35 325
rect -15 55 0 325
rect -50 40 0 55
rect 50 325 100 340
rect 50 55 65 325
rect 85 55 100 325
rect 50 40 100 55
rect 150 325 200 340
rect 150 55 165 325
rect 185 55 200 325
rect 150 40 200 55
rect 230 325 280 340
rect 230 55 245 325
rect 265 55 280 325
rect 230 40 280 55
rect 330 325 380 340
rect 330 55 345 325
rect 365 55 380 325
rect 330 40 380 55
rect 430 325 480 340
rect 430 55 445 325
rect 465 55 480 325
rect 430 40 480 55
rect 510 325 560 340
rect 510 55 525 325
rect 545 55 560 325
rect 510 40 560 55
rect 610 325 660 340
rect 610 55 625 325
rect 645 55 660 325
rect 610 40 660 55
rect 710 325 760 340
rect 710 55 725 325
rect 745 55 760 325
rect 710 40 760 55
rect 790 325 840 340
rect 790 55 805 325
rect 825 55 840 325
rect 790 40 840 55
rect 890 325 940 340
rect 890 55 905 325
rect 925 55 940 325
rect 890 40 940 55
rect 990 325 1040 340
rect 990 55 1005 325
rect 1025 55 1040 325
rect 990 40 1040 55
rect 1070 325 1120 340
rect 1070 55 1085 325
rect 1105 55 1120 325
rect 1070 40 1120 55
rect 1170 325 1220 340
rect 1170 55 1185 325
rect 1205 55 1220 325
rect 1170 40 1220 55
rect 1270 325 1320 340
rect 1270 55 1285 325
rect 1305 55 1320 325
rect 1270 40 1320 55
rect 110 -85 160 -70
rect 110 -355 125 -85
rect 145 -355 160 -85
rect 110 -370 160 -355
rect 210 -85 260 -70
rect 210 -355 225 -85
rect 245 -355 260 -85
rect 210 -370 260 -355
rect 310 -85 360 -70
rect 310 -355 325 -85
rect 345 -355 360 -85
rect 310 -370 360 -355
rect 410 -85 460 -70
rect 410 -355 425 -85
rect 445 -355 460 -85
rect 410 -370 460 -355
rect 510 -85 560 -70
rect 510 -355 525 -85
rect 545 -355 560 -85
rect 510 -370 560 -355
rect 610 -85 660 -70
rect 610 -355 625 -85
rect 645 -355 660 -85
rect 610 -370 660 -355
rect 710 -85 760 -70
rect 710 -355 725 -85
rect 745 -355 760 -85
rect 710 -370 760 -355
rect 810 -85 860 -70
rect 810 -355 825 -85
rect 845 -355 860 -85
rect 810 -370 860 -355
rect 910 -85 960 -70
rect 910 -355 925 -85
rect 945 -355 960 -85
rect 910 -370 960 -355
rect 1010 -85 1060 -70
rect 1010 -355 1025 -85
rect 1045 -355 1060 -85
rect 1010 -370 1060 -355
rect 1110 -85 1160 -70
rect 1110 -355 1125 -85
rect 1145 -355 1160 -85
rect 1110 -370 1160 -355
<< pdiff >>
rect 110 2125 160 2140
rect 110 1355 125 2125
rect 145 1355 160 2125
rect 110 1340 160 1355
rect 210 2125 260 2140
rect 210 1355 225 2125
rect 245 1355 260 2125
rect 210 1340 260 1355
rect 310 2125 360 2140
rect 310 1355 325 2125
rect 345 1355 360 2125
rect 310 1340 360 1355
rect 410 2125 460 2140
rect 410 1355 425 2125
rect 445 1355 460 2125
rect 410 1340 460 1355
rect 510 2125 560 2140
rect 510 1355 525 2125
rect 545 1355 560 2125
rect 510 1340 560 1355
rect 610 2125 660 2140
rect 610 1355 625 2125
rect 645 1355 660 2125
rect 610 1340 660 1355
rect 710 2125 760 2140
rect 710 1355 725 2125
rect 745 1355 760 2125
rect 710 1340 760 1355
rect 810 2125 860 2140
rect 810 1355 825 2125
rect 845 1355 860 2125
rect 810 1340 860 1355
rect 910 2125 960 2140
rect 910 1355 925 2125
rect 945 1355 960 2125
rect 910 1340 960 1355
rect 1010 2125 1060 2140
rect 1010 1355 1025 2125
rect 1045 1355 1060 2125
rect 1010 1340 1060 1355
rect 1110 2125 1160 2140
rect 1110 1355 1125 2125
rect 1145 1355 1160 2125
rect 1110 1340 1160 1355
rect -50 1180 0 1195
rect -50 410 -35 1180
rect -15 410 0 1180
rect -50 395 0 410
rect 50 1180 100 1195
rect 50 410 65 1180
rect 85 410 100 1180
rect 50 395 100 410
rect 150 1180 200 1195
rect 150 410 165 1180
rect 185 410 200 1180
rect 150 395 200 410
rect 230 1180 280 1195
rect 230 410 245 1180
rect 265 410 280 1180
rect 230 395 280 410
rect 330 1180 380 1195
rect 330 410 345 1180
rect 365 410 380 1180
rect 330 395 380 410
rect 430 1180 480 1195
rect 430 410 445 1180
rect 465 410 480 1180
rect 430 395 480 410
rect 510 1180 560 1195
rect 510 410 525 1180
rect 545 410 560 1180
rect 510 395 560 410
rect 610 1180 660 1195
rect 610 410 625 1180
rect 645 410 660 1180
rect 610 395 660 410
rect 710 1180 760 1195
rect 710 410 725 1180
rect 745 410 760 1180
rect 710 395 760 410
rect 790 1180 840 1195
rect 790 410 805 1180
rect 825 410 840 1180
rect 790 395 840 410
rect 890 1180 940 1195
rect 890 410 905 1180
rect 925 410 940 1180
rect 890 395 940 410
rect 990 1180 1040 1195
rect 990 410 1005 1180
rect 1025 410 1040 1180
rect 990 395 1040 410
rect 1070 1180 1120 1195
rect 1070 410 1085 1180
rect 1105 410 1120 1180
rect 1070 395 1120 410
rect 1170 1180 1220 1195
rect 1170 410 1185 1180
rect 1205 410 1220 1180
rect 1170 395 1220 410
rect 1270 1180 1320 1195
rect 1270 410 1285 1180
rect 1305 410 1320 1180
rect 1270 395 1320 410
<< ndiffc >>
rect -35 55 -15 325
rect 65 55 85 325
rect 165 55 185 325
rect 245 55 265 325
rect 345 55 365 325
rect 445 55 465 325
rect 525 55 545 325
rect 625 55 645 325
rect 725 55 745 325
rect 805 55 825 325
rect 905 55 925 325
rect 1005 55 1025 325
rect 1085 55 1105 325
rect 1185 55 1205 325
rect 1285 55 1305 325
rect 125 -355 145 -85
rect 225 -355 245 -85
rect 325 -355 345 -85
rect 425 -355 445 -85
rect 525 -355 545 -85
rect 625 -355 645 -85
rect 725 -355 745 -85
rect 825 -355 845 -85
rect 925 -355 945 -85
rect 1025 -355 1045 -85
rect 1125 -355 1145 -85
<< pdiffc >>
rect 125 1355 145 2125
rect 225 1355 245 2125
rect 325 1355 345 2125
rect 425 1355 445 2125
rect 525 1355 545 2125
rect 625 1355 645 2125
rect 725 1355 745 2125
rect 825 1355 845 2125
rect 925 1355 945 2125
rect 1025 1355 1045 2125
rect 1125 1355 1145 2125
rect -35 410 -15 1180
rect 65 410 85 1180
rect 165 410 185 1180
rect 245 410 265 1180
rect 345 410 365 1180
rect 445 410 465 1180
rect 525 410 545 1180
rect 625 410 645 1180
rect 725 410 745 1180
rect 805 410 825 1180
rect 905 410 925 1180
rect 1005 410 1025 1180
rect 1085 410 1105 1180
rect 1185 410 1205 1180
rect 1285 410 1305 1180
<< psubdiff >>
rect -50 -85 110 -70
rect -50 -355 -35 -85
rect 100 -355 110 -85
rect -50 -370 110 -355
rect 1160 -85 1320 -70
rect 1160 -355 1170 -85
rect 1305 -355 1320 -85
rect 1160 -370 1320 -355
<< nsubdiff >>
rect -50 2125 110 2140
rect -50 1355 -35 2125
rect 95 1355 110 2125
rect -50 1340 110 1355
rect 1160 2125 1320 2140
rect 1160 1355 1175 2125
rect 1305 1355 1320 2125
rect 1160 1340 1320 1355
<< psubdiffcont >>
rect -35 -355 100 -85
rect 1170 -355 1305 -85
<< nsubdiffcont >>
rect -35 1355 95 2125
rect 1175 1355 1305 2125
<< poly >>
rect 165 2215 310 2230
rect 165 2195 175 2215
rect 195 2205 310 2215
rect 195 2195 1010 2205
rect 165 2180 1010 2195
rect 260 2155 1010 2180
rect 160 2140 210 2155
rect 260 2140 310 2155
rect 360 2140 410 2155
rect 460 2140 510 2155
rect 560 2140 610 2155
rect 660 2140 710 2155
rect 760 2140 810 2155
rect 860 2140 910 2155
rect 960 2140 1010 2155
rect 1060 2140 1110 2155
rect 55 1310 125 1325
rect 55 1290 65 1310
rect 85 1290 125 1310
rect 55 1275 125 1290
rect 160 1315 210 1340
rect 260 1325 310 1340
rect 360 1325 410 1340
rect 460 1325 510 1340
rect 560 1325 610 1340
rect 660 1325 710 1340
rect 760 1325 810 1340
rect 860 1325 910 1340
rect 960 1325 1010 1340
rect 160 1295 175 1315
rect 195 1295 210 1315
rect 160 1285 210 1295
rect 1060 1315 1110 1340
rect 1060 1295 1075 1315
rect 1095 1295 1110 1315
rect 1060 1285 1110 1295
rect 75 1260 125 1275
rect 0 1240 50 1250
rect 0 1220 15 1240
rect 35 1220 50 1240
rect 0 1195 50 1220
rect 75 1210 1170 1260
rect 100 1195 150 1210
rect 280 1195 330 1210
rect 380 1195 430 1210
rect 560 1195 610 1210
rect 660 1195 710 1210
rect 840 1195 890 1210
rect 940 1195 990 1210
rect 1120 1195 1170 1210
rect 1220 1240 1270 1250
rect 1220 1220 1235 1240
rect 1255 1220 1270 1240
rect 1220 1195 1270 1220
rect 0 380 50 395
rect 100 380 150 395
rect 280 380 330 395
rect 380 380 430 395
rect 560 380 610 395
rect 660 380 710 395
rect 840 380 890 395
rect 940 380 990 395
rect 1120 380 1170 395
rect 1220 380 1270 395
rect 0 340 50 355
rect 100 340 150 355
rect 280 340 330 355
rect 380 340 430 355
rect 560 340 610 355
rect 660 340 710 355
rect 840 340 890 355
rect 940 340 990 355
rect 1120 340 1170 355
rect 1220 340 1270 355
rect 0 15 50 40
rect 100 25 150 40
rect 280 25 330 40
rect 380 25 430 40
rect 560 25 610 40
rect 660 25 710 40
rect 840 25 890 40
rect 940 25 990 40
rect 1120 25 1170 40
rect 0 -5 15 15
rect 35 -5 50 15
rect 0 -15 50 -5
rect 85 -25 1170 25
rect 1220 15 1270 40
rect 1220 -5 1235 15
rect 1255 -5 1270 15
rect 1220 -15 1270 -5
rect 85 -45 100 -25
rect 120 -45 135 -25
rect 85 -55 135 -45
rect 160 -70 210 -55
rect 260 -70 310 -55
rect 360 -70 410 -55
rect 460 -70 510 -55
rect 560 -70 610 -55
rect 660 -70 710 -55
rect 760 -70 810 -55
rect 860 -70 910 -55
rect 960 -70 1010 -55
rect 1060 -70 1110 -55
rect 160 -395 210 -370
rect 160 -415 175 -395
rect 195 -415 210 -395
rect 160 -425 210 -415
rect 260 -385 310 -370
rect 360 -385 410 -370
rect 460 -385 510 -370
rect 560 -385 610 -370
rect 660 -385 710 -370
rect 760 -385 810 -370
rect 860 -385 910 -370
rect 960 -385 1010 -370
rect 260 -395 1010 -385
rect 260 -415 575 -395
rect 595 -415 675 -395
rect 695 -415 1010 -395
rect 260 -435 1010 -415
rect 1060 -395 1110 -370
rect 1060 -415 1075 -395
rect 1095 -415 1110 -395
rect 1060 -425 1110 -415
<< polycont >>
rect 175 2195 195 2215
rect 65 1290 85 1310
rect 175 1295 195 1315
rect 1075 1295 1095 1315
rect 15 1220 35 1240
rect 1235 1220 1255 1240
rect 15 -5 35 15
rect 1235 -5 1255 15
rect 100 -45 120 -25
rect 175 -415 195 -395
rect 575 -415 595 -395
rect 675 -415 695 -395
rect 1075 -415 1095 -395
<< locali >>
rect 225 2230 1045 2250
rect 165 2215 205 2225
rect 165 2205 175 2215
rect -50 2195 175 2205
rect 195 2195 205 2215
rect -50 2185 205 2195
rect 225 2210 245 2230
rect 225 2200 265 2210
rect 225 2180 235 2200
rect 255 2180 265 2200
rect 225 2170 265 2180
rect 415 2200 455 2210
rect 415 2180 425 2200
rect 445 2180 455 2200
rect 415 2170 455 2180
rect 225 2135 245 2170
rect 425 2135 445 2170
rect 625 2135 645 2230
rect 815 2200 855 2210
rect 815 2180 825 2200
rect 845 2180 855 2200
rect 815 2170 855 2180
rect 825 2135 845 2170
rect 1025 2135 1045 2230
rect -45 2125 155 2135
rect -45 1355 -35 2125
rect 95 1355 125 2125
rect 145 1355 155 2125
rect -45 1345 155 1355
rect 215 2125 255 2135
rect 215 1355 225 2125
rect 245 1355 255 2125
rect 215 1345 255 1355
rect 315 2125 355 2135
rect 315 1355 325 2125
rect 345 1355 355 2125
rect 315 1345 355 1355
rect 415 2125 455 2135
rect 415 1355 425 2125
rect 445 1355 455 2125
rect 415 1345 455 1355
rect 515 2125 555 2135
rect 515 1355 525 2125
rect 545 1355 555 2125
rect 515 1345 555 1355
rect 615 2125 655 2135
rect 615 1355 625 2125
rect 645 1355 655 2125
rect 615 1345 655 1355
rect 715 2125 755 2135
rect 715 1355 725 2125
rect 745 1355 755 2125
rect 715 1345 755 1355
rect 815 2125 855 2135
rect 815 1355 825 2125
rect 845 1355 855 2125
rect 815 1345 855 1355
rect 915 2125 955 2135
rect 915 1355 925 2125
rect 945 1355 955 2125
rect 915 1345 955 1355
rect 1015 2125 1055 2135
rect 1015 1355 1025 2125
rect 1045 1355 1055 2125
rect 1015 1345 1055 1355
rect 1115 2125 1315 2135
rect 1115 1355 1125 2125
rect 1145 1355 1175 2125
rect 1305 1355 1315 2125
rect 1115 1345 1315 1355
rect 115 1325 155 1345
rect 55 1310 95 1320
rect 55 1300 65 1310
rect -50 1290 65 1300
rect 85 1290 95 1310
rect -50 1280 95 1290
rect 115 1315 205 1325
rect 115 1295 175 1315
rect 195 1295 205 1315
rect 115 1285 205 1295
rect -45 1240 45 1250
rect -45 1220 15 1240
rect 35 1220 45 1240
rect 225 1230 245 1345
rect 425 1230 445 1345
rect -45 1210 45 1220
rect 65 1210 245 1230
rect 345 1210 445 1230
rect -45 1180 -5 1210
rect 65 1190 85 1210
rect 345 1190 365 1210
rect 625 1190 645 1345
rect 825 1230 845 1345
rect 1025 1230 1045 1345
rect 1115 1325 1155 1345
rect 1065 1315 1155 1325
rect 1065 1295 1075 1315
rect 1095 1295 1155 1315
rect 1065 1285 1155 1295
rect 1225 1240 1315 1250
rect 825 1210 925 1230
rect 1025 1210 1205 1230
rect 1225 1220 1235 1240
rect 1255 1220 1315 1240
rect 1225 1210 1315 1220
rect 905 1190 925 1210
rect 1185 1190 1205 1210
rect -45 410 -35 1180
rect -15 410 -5 1180
rect -45 400 -5 410
rect 55 1180 95 1190
rect 55 410 65 1180
rect 85 410 95 1180
rect 55 400 95 410
rect 155 1180 195 1190
rect 155 410 165 1180
rect 185 410 195 1180
rect 155 400 195 410
rect 235 1180 275 1190
rect 235 410 245 1180
rect 265 410 275 1180
rect 235 400 275 410
rect 335 1180 375 1190
rect 335 410 345 1180
rect 365 410 375 1180
rect 335 400 375 410
rect 435 1180 475 1190
rect 435 410 445 1180
rect 465 410 475 1180
rect 435 400 475 410
rect 515 1180 555 1190
rect 515 410 525 1180
rect 545 410 555 1180
rect 515 400 555 410
rect 615 1180 655 1190
rect 615 410 625 1180
rect 645 410 655 1180
rect 615 400 655 410
rect 715 1180 755 1190
rect 715 410 725 1180
rect 745 410 755 1180
rect 715 400 755 410
rect 795 1180 835 1190
rect 795 410 805 1180
rect 825 410 835 1180
rect 795 400 835 410
rect 895 1180 935 1190
rect 895 410 905 1180
rect 925 410 935 1180
rect 895 400 935 410
rect 995 1180 1035 1190
rect 995 410 1005 1180
rect 1025 410 1035 1180
rect 995 400 1035 410
rect 1075 1180 1115 1190
rect 1075 410 1085 1180
rect 1105 410 1115 1180
rect 1075 400 1115 410
rect 1175 1180 1215 1190
rect 1175 410 1185 1180
rect 1205 410 1215 1180
rect 1175 400 1215 410
rect 1275 1180 1315 1210
rect 1275 410 1285 1180
rect 1305 410 1315 1180
rect 1275 400 1315 410
rect 165 335 185 400
rect 245 335 265 400
rect 445 335 465 400
rect 525 335 545 400
rect 725 335 745 400
rect 805 335 825 400
rect 1005 335 1025 400
rect 1085 335 1105 400
rect -45 325 -5 335
rect -45 55 -35 325
rect -15 55 -5 325
rect -45 25 -5 55
rect 55 325 95 335
rect 55 55 65 325
rect 85 65 95 325
rect 155 325 195 335
rect 85 55 135 65
rect 55 45 135 55
rect 155 55 165 325
rect 185 55 195 325
rect 155 45 195 55
rect 235 325 275 335
rect 235 55 245 325
rect 265 55 275 325
rect 235 45 275 55
rect 335 325 375 335
rect 335 55 345 325
rect 365 55 375 325
rect 335 45 375 55
rect 435 325 475 335
rect 435 55 445 325
rect 465 55 475 325
rect 435 45 475 55
rect 515 325 555 335
rect 515 55 525 325
rect 545 55 555 325
rect 515 45 555 55
rect 615 325 655 335
rect 615 55 625 325
rect 645 55 655 325
rect 615 45 655 55
rect 715 325 755 335
rect 715 55 725 325
rect 745 55 755 325
rect 715 45 755 55
rect 795 325 835 335
rect 795 55 805 325
rect 825 55 835 325
rect 795 45 835 55
rect 895 325 935 335
rect 895 55 905 325
rect 925 55 935 325
rect 895 45 935 55
rect 995 325 1035 335
rect 995 55 1005 325
rect 1025 55 1035 325
rect 995 45 1035 55
rect 1075 325 1115 335
rect 1075 55 1085 325
rect 1105 55 1115 325
rect 1075 45 1115 55
rect 1175 325 1215 335
rect 1175 55 1185 325
rect 1205 55 1215 325
rect 1175 45 1215 55
rect 1275 325 1315 335
rect 1275 55 1285 325
rect 1305 55 1315 325
rect 115 25 135 45
rect 345 25 365 45
rect 525 25 545 45
rect -45 15 45 25
rect -45 -5 15 15
rect 35 -5 45 15
rect 115 5 245 25
rect 345 5 445 25
rect 525 5 595 25
rect -45 -15 45 -5
rect 90 -25 130 -15
rect 90 -35 100 -25
rect -50 -45 100 -35
rect 120 -45 130 -25
rect -50 -55 130 -45
rect 225 -75 245 5
rect 425 -75 445 5
rect -45 -85 155 -75
rect -45 -355 -35 -85
rect 100 -355 125 -85
rect 145 -355 155 -85
rect -45 -365 155 -355
rect 215 -85 255 -75
rect 215 -355 225 -85
rect 245 -355 255 -85
rect 215 -365 255 -355
rect 315 -85 355 -75
rect 315 -355 325 -85
rect 345 -355 355 -85
rect 315 -365 355 -355
rect 415 -85 455 -75
rect 415 -355 425 -85
rect 445 -355 455 -85
rect 415 -365 455 -355
rect 515 -85 555 -75
rect 515 -355 525 -85
rect 545 -355 555 -85
rect 515 -365 555 -355
rect 115 -385 155 -365
rect 575 -385 595 5
rect 625 -75 645 45
rect 725 25 745 45
rect 905 25 925 45
rect 1185 25 1205 45
rect 1275 25 1315 55
rect 675 5 745 25
rect 825 5 925 25
rect 1025 5 1205 25
rect 1225 15 1315 25
rect 615 -85 655 -75
rect 615 -355 625 -85
rect 645 -355 655 -85
rect 615 -365 655 -355
rect 675 -385 695 5
rect 825 -75 845 5
rect 1025 -75 1045 5
rect 1225 -5 1235 15
rect 1255 -5 1315 15
rect 1225 -15 1315 -5
rect 715 -85 755 -75
rect 715 -355 725 -85
rect 745 -355 755 -85
rect 715 -365 755 -355
rect 815 -85 855 -75
rect 815 -355 825 -85
rect 845 -355 855 -85
rect 815 -365 855 -355
rect 915 -85 955 -75
rect 915 -355 925 -85
rect 945 -355 955 -85
rect 915 -365 955 -355
rect 1015 -85 1055 -75
rect 1015 -355 1025 -85
rect 1045 -355 1055 -85
rect 1015 -365 1055 -355
rect 1115 -85 1315 -75
rect 1115 -355 1125 -85
rect 1145 -355 1170 -85
rect 1305 -355 1315 -85
rect 1115 -365 1315 -355
rect 1115 -385 1155 -365
rect 115 -395 205 -385
rect 115 -415 175 -395
rect 195 -415 205 -395
rect 115 -425 205 -415
rect 565 -395 605 -385
rect 565 -415 575 -395
rect 595 -415 605 -395
rect 565 -425 605 -415
rect 665 -395 705 -385
rect 665 -415 675 -395
rect 695 -415 705 -395
rect 665 -425 705 -415
rect 1065 -395 1155 -385
rect 1065 -415 1075 -395
rect 1095 -415 1155 -395
rect 1065 -425 1155 -415
<< viali >>
rect 235 2180 255 2200
rect 425 2180 445 2200
rect 825 2180 845 2200
rect -35 1355 95 2125
rect 125 1355 145 2125
rect 325 1355 345 2125
rect 525 1355 545 2125
rect 725 1355 745 2125
rect 925 1355 945 2125
rect 1125 1355 1145 2125
rect 1175 1355 1305 2125
rect 15 1220 35 1240
rect 1235 1220 1255 1240
rect 65 410 85 430
rect 345 440 365 460
rect 625 410 645 430
rect 905 440 925 460
rect 1185 410 1205 430
rect 65 305 85 325
rect 165 245 185 265
rect 245 190 265 210
rect 345 275 365 295
rect 445 190 465 210
rect 525 220 545 240
rect 625 305 645 325
rect 725 220 745 240
rect 805 190 825 210
rect 905 275 925 295
rect 1005 190 1025 210
rect 1085 245 1105 265
rect 1185 305 1205 325
rect 15 -5 35 15
rect -35 -355 100 -85
rect 125 -355 145 -85
rect 325 -355 345 -85
rect 525 -355 545 -85
rect 1235 -5 1255 15
rect 725 -355 745 -85
rect 925 -355 945 -85
rect 1125 -355 1145 -85
rect 1170 -355 1305 -85
<< metal1 >>
rect 235 2210 265 2250
rect 225 2200 265 2210
rect 225 2180 235 2200
rect 255 2180 265 2200
rect 225 2170 265 2180
rect 415 2210 445 2250
rect 415 2200 455 2210
rect 815 2200 855 2210
rect 415 2180 425 2200
rect 445 2180 825 2200
rect 845 2180 855 2200
rect 415 2170 855 2180
rect -50 2125 1320 2140
rect -50 1355 -35 2125
rect 95 1355 125 2125
rect 145 1355 325 2125
rect 345 1355 525 2125
rect 545 1355 725 2125
rect 745 1355 925 2125
rect 945 1355 1125 2125
rect 1145 1355 1175 2125
rect 1305 1355 1320 2125
rect -50 1340 1320 1355
rect 5 1240 45 1340
rect 5 1220 15 1240
rect 35 1220 45 1240
rect 5 1210 45 1220
rect 1225 1240 1265 1340
rect 1225 1220 1235 1240
rect 1255 1220 1265 1240
rect 1225 1210 1265 1220
rect 335 460 935 470
rect 335 440 345 460
rect 365 455 905 460
rect 365 440 375 455
rect 895 440 905 455
rect 925 440 935 460
rect 55 430 95 440
rect 335 430 375 440
rect 615 430 655 440
rect 895 430 935 440
rect 1175 430 1215 440
rect 55 410 65 430
rect 85 415 95 430
rect 615 415 625 430
rect 85 410 625 415
rect 645 415 655 430
rect 1175 415 1185 430
rect 645 410 1185 415
rect 1205 410 1215 430
rect 55 400 1215 410
rect 55 325 1215 335
rect 55 305 65 325
rect 85 320 625 325
rect 85 305 95 320
rect 615 305 625 320
rect 645 320 1185 325
rect 645 305 655 320
rect 1175 305 1185 320
rect 1205 305 1215 325
rect 55 295 95 305
rect 335 295 375 305
rect 615 295 655 305
rect 895 295 935 305
rect 1175 295 1215 305
rect 335 275 345 295
rect 365 280 375 295
rect 895 280 905 295
rect 365 275 905 280
rect 925 275 935 295
rect 155 265 195 275
rect 335 265 935 275
rect 1075 265 1115 275
rect 155 245 165 265
rect 185 250 195 265
rect 1075 250 1085 265
rect 185 245 1085 250
rect 1105 245 1115 265
rect 155 240 1115 245
rect 155 235 525 240
rect 515 220 525 235
rect 545 235 725 240
rect 545 220 555 235
rect 235 210 275 220
rect 235 190 245 210
rect 265 195 275 210
rect 435 210 475 220
rect 515 210 555 220
rect 715 220 725 235
rect 745 235 1115 240
rect 745 220 755 235
rect 715 210 755 220
rect 795 210 835 220
rect 435 195 445 210
rect 265 190 445 195
rect 465 195 475 210
rect 795 195 805 210
rect 465 190 805 195
rect 825 195 835 210
rect 995 210 1035 220
rect 995 195 1005 210
rect 825 190 1005 195
rect 1025 195 1035 210
rect 1025 190 1410 195
rect 235 180 1410 190
rect 5 15 45 25
rect 5 -5 15 15
rect 35 -5 45 15
rect 5 -70 45 -5
rect 1225 15 1265 25
rect 1225 -5 1235 15
rect 1255 -5 1265 15
rect 1225 -70 1265 -5
rect -50 -85 1320 -70
rect -50 -355 -35 -85
rect 100 -355 125 -85
rect 145 -355 325 -85
rect 345 -355 525 -85
rect 545 -355 725 -85
rect 745 -355 925 -85
rect 945 -355 1125 -85
rect 1145 -355 1170 -85
rect 1305 -355 1320 -85
rect -50 -370 1320 -355
<< labels >>
flabel metal1 1410 190 1410 190 3 FreeSans 160 0 0 0 Vout
port 3 e
flabel locali -50 -45 -50 -45 7 FreeSans 160 0 0 0 Vcn
port 5 w
flabel metal1 -50 -220 -50 -220 7 FreeSans 160 0 0 0 VN
port 9 w
flabel locali -50 1290 -50 1290 7 FreeSans 160 0 0 0 Vcp
port 6 w
flabel metal1 -50 1490 -50 1490 7 FreeSans 160 0 0 0 VP
port 8 w
flabel locali -50 2195 -50 2195 7 FreeSans 160 0 0 0 Vbp
port 7 w
flabel metal1 250 2250 250 2250 1 FreeSans 160 0 0 0 I1
port 1 n
flabel metal1 430 2250 430 2250 1 FreeSans 160 0 0 0 I2
port 2 n
<< end >>
