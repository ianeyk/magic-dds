magic
tech sky130A
timestamp 1702426134
<< error_s >>
rect 0 6535 17 6547
rect -17 6520 0 6530
rect -10 6518 0 6520
rect -135 5300 -133 5310
rect -152 5290 -150 5300
<< locali >>
rect -3580 1395 -3560 8225
rect -3540 2710 -3520 8225
rect -3500 4025 -3480 8225
rect -3460 5340 -3440 8225
rect -2520 8215 -2480 8225
rect -2520 8195 -2510 8215
rect -2490 8195 -2480 8215
rect -2520 8100 -2480 8195
rect -2520 8080 -2510 8100
rect -2490 8080 -2480 8100
rect -2520 8070 -2480 8080
rect -2090 7970 -2070 8225
rect -2050 8030 -2030 8225
rect -2010 8070 -1990 8225
rect -1970 8110 -1950 8225
rect -1870 8215 -1830 8225
rect -1870 8195 -1860 8215
rect -1840 8195 -1830 8215
rect -1970 8090 -1930 8110
rect -2010 8050 -1970 8070
rect -2050 8020 -2010 8030
rect -2050 8000 -2040 8020
rect -2020 8000 -2010 8020
rect -2050 7990 -2010 8000
rect -1990 8010 -1970 8050
rect -1950 8050 -1930 8090
rect -1870 8100 -1830 8195
rect -1220 8215 -1180 8225
rect -1220 8195 -1210 8215
rect -1190 8195 -1180 8215
rect -1870 8080 -1860 8100
rect -1840 8080 -1830 8100
rect -1870 8070 -1830 8080
rect -1560 8090 -1320 8110
rect -1560 8050 -1540 8090
rect -1400 8060 -1360 8070
rect -1400 8050 -1390 8060
rect -1950 8030 -1540 8050
rect -1520 8040 -1390 8050
rect -1370 8040 -1360 8060
rect -1520 8030 -1360 8040
rect -1340 8050 -1320 8090
rect -1220 8100 -1180 8195
rect -570 8215 -530 8225
rect -570 8195 -560 8215
rect -540 8195 -530 8215
rect -1220 8080 -1210 8100
rect -1190 8080 -1180 8100
rect -1220 8070 -1180 8080
rect -910 8100 -710 8110
rect -910 8090 -740 8100
rect -910 8050 -890 8090
rect -750 8080 -740 8090
rect -720 8080 -710 8100
rect -750 8070 -710 8080
rect -570 8100 -530 8195
rect -570 8080 -560 8100
rect -540 8080 -530 8100
rect -570 8070 -530 8080
rect 1030 8215 1070 8225
rect 1030 8195 1040 8215
rect 1060 8195 1070 8215
rect 1030 8100 1070 8195
rect 1030 8080 1040 8100
rect 1060 8080 1070 8100
rect 1030 8070 1070 8080
rect 1680 8215 1720 8225
rect 1680 8195 1690 8215
rect 1710 8195 1720 8215
rect 1680 8100 1720 8195
rect 1680 8080 1690 8100
rect 1710 8080 1720 8100
rect 1680 8070 1720 8080
rect 2330 8215 2370 8225
rect 2330 8195 2340 8215
rect 2360 8195 2370 8215
rect 2330 8100 2370 8195
rect 2330 8080 2340 8100
rect 2360 8080 2370 8100
rect 2330 8070 2370 8080
rect 2980 8215 3020 8225
rect 2980 8195 2990 8215
rect 3010 8195 3020 8215
rect 2980 8100 3020 8195
rect 2980 8080 2990 8100
rect 3010 8080 3020 8100
rect 2980 8070 3020 8080
rect -1340 8030 -890 8050
rect -870 8030 140 8050
rect -1520 8010 -1500 8030
rect -870 8010 -850 8030
rect 120 8010 140 8030
rect -1990 7990 -1500 8010
rect -1480 7990 -850 8010
rect -830 7990 100 8010
rect 120 7990 710 8010
rect -1480 7970 -1460 7990
rect -830 7970 -810 7990
rect 80 7970 100 7990
rect 690 7970 710 7990
rect -2090 7950 -1460 7970
rect -1440 7950 -810 7970
rect -790 7950 60 7970
rect 80 7950 670 7970
rect 690 7950 1320 7970
rect -2090 7930 -2070 7950
rect -1440 7930 -1420 7950
rect -790 7930 -770 7950
rect 40 7930 60 7950
rect 650 7930 670 7950
rect 1300 7930 1320 7950
rect -3420 7920 -3380 7930
rect -3420 7900 -3410 7920
rect -3390 7900 -3380 7920
rect -3420 7890 -3380 7900
rect -3350 7920 -3310 7930
rect -3350 7900 -3340 7920
rect -3320 7900 -3310 7920
rect -3350 7890 -3310 7900
rect -2700 7920 -2070 7930
rect -2700 7900 -2690 7920
rect -2670 7910 -2070 7920
rect -2050 7920 -1420 7930
rect -2670 7900 -2660 7910
rect -2700 7890 -2660 7900
rect -2050 7900 -2040 7920
rect -2020 7910 -1420 7920
rect -1400 7920 -770 7930
rect -2020 7900 -2010 7910
rect -2050 7890 -2010 7900
rect -1400 7900 -1390 7920
rect -1370 7910 -770 7920
rect -750 7920 0 7930
rect -1370 7900 -1360 7910
rect -1400 7890 -1360 7900
rect -750 7900 -740 7920
rect -720 7910 0 7920
rect 40 7910 630 7930
rect 650 7910 1280 7930
rect 1300 7910 1930 7930
rect -720 7900 -710 7910
rect -750 7890 -710 7900
rect -3420 6655 -3400 7890
rect -20 7850 0 7910
rect 610 7890 630 7910
rect 1260 7890 1280 7910
rect 1910 7890 1930 7910
rect -130 7810 0 7830
rect -130 6655 -110 7810
rect -3420 6635 -3380 6655
rect -150 6635 -110 6655
rect -40 6520 0 6530
rect -40 6500 -30 6520
rect -10 6500 0 6520
rect -40 6490 0 6500
rect -3460 5320 -3380 5340
rect -150 5330 -95 5340
rect -150 5320 -125 5330
rect -135 5310 -125 5320
rect -105 5310 -95 5330
rect -135 5300 -95 5310
rect -135 5190 0 5200
rect -135 5170 -125 5190
rect -105 5180 0 5190
rect -105 5170 -95 5180
rect -135 5160 -95 5170
rect -3500 4005 -3380 4025
rect -150 4005 -110 4025
rect -130 3885 -110 4005
rect -130 3865 0 3885
rect -135 2720 -95 2730
rect -135 2710 -125 2720
rect -3540 2690 -3380 2710
rect -150 2700 -125 2710
rect -105 2700 -95 2720
rect -150 2690 -95 2700
rect -95 2580 -55 2590
rect -95 2560 -85 2580
rect -65 2570 -55 2580
rect -65 2560 0 2570
rect -95 2550 0 2560
rect -65 1405 -25 1415
rect -65 1395 -55 1405
rect -3580 1375 -3380 1395
rect -150 1385 -55 1395
rect -35 1385 -25 1405
rect -150 1375 -25 1385
rect -130 1235 0 1255
rect -130 80 -110 1235
rect -3470 70 -3380 80
rect -3470 50 -3460 70
rect -3440 60 -3380 70
rect -150 60 -110 80
rect -3440 50 -3430 60
rect -3470 40 -3430 50
rect -3280 -10 -3240 0
rect -3280 -30 -3270 -10
rect -3250 -30 -3240 -10
rect -3280 -140 -3240 -30
rect -3280 -160 -3270 -140
rect -3250 -160 -3240 -140
rect -3280 -170 -3240 -160
rect -2630 -10 -2590 0
rect -2630 -30 -2620 -10
rect -2600 -30 -2590 -10
rect -2630 -140 -2590 -30
rect -2630 -160 -2620 -140
rect -2600 -160 -2590 -140
rect -2630 -170 -2590 -160
rect -1980 -10 -1940 0
rect -1980 -30 -1970 -10
rect -1950 -30 -1940 -10
rect -1980 -140 -1940 -30
rect -1980 -160 -1970 -140
rect -1950 -160 -1940 -140
rect -1980 -170 -1940 -160
rect -1330 -10 -1290 0
rect -1330 -30 -1320 -10
rect -1300 -30 -1290 -10
rect -1330 -140 -1290 -30
rect -1330 -160 -1320 -140
rect -1300 -160 -1290 -140
rect -1330 -170 -1290 -160
rect -680 -10 -640 0
rect -680 -30 -670 -10
rect -650 -30 -640 -10
rect -680 -140 -640 -30
rect -680 -160 -670 -140
rect -650 -160 -640 -140
rect -680 -170 -640 -160
rect 505 -10 545 0
rect 505 -30 515 -10
rect 535 -30 545 -10
rect 505 -140 545 -30
rect 505 -160 515 -140
rect 535 -160 545 -140
rect 505 -170 545 -160
rect 1155 -10 1195 0
rect 1155 -30 1165 -10
rect 1185 -30 1195 -10
rect 1155 -140 1195 -30
rect 1155 -160 1165 -140
rect 1185 -160 1195 -140
rect 1155 -170 1195 -160
rect 1805 -10 1845 0
rect 1805 -30 1815 -10
rect 1835 -30 1845 -10
rect 1805 -140 1845 -30
rect 1805 -160 1815 -140
rect 1835 -160 1845 -140
rect 1805 -170 1845 -160
rect 2455 -10 2495 0
rect 2455 -30 2465 -10
rect 2485 -30 2495 -10
rect 2455 -140 2495 -30
rect 2455 -160 2465 -140
rect 2485 -160 2495 -140
rect 2455 -170 2495 -160
rect 3105 -10 3145 0
rect 3105 -30 3115 -10
rect 3135 -30 3145 -10
rect 3105 -140 3145 -30
rect 3105 -160 3115 -140
rect 3135 -160 3145 -140
rect 3105 -170 3145 -160
<< viali >>
rect -2510 8195 -2490 8215
rect -2510 8080 -2490 8100
rect -1860 8195 -1840 8215
rect -2040 8000 -2020 8020
rect -1210 8195 -1190 8215
rect -1860 8080 -1840 8100
rect -1390 8040 -1370 8060
rect -560 8195 -540 8215
rect -1210 8080 -1190 8100
rect -740 8080 -720 8100
rect -560 8080 -540 8100
rect 1040 8195 1060 8215
rect 1040 8080 1060 8100
rect 1690 8195 1710 8215
rect 1690 8080 1710 8100
rect 2340 8195 2360 8215
rect 2340 8080 2360 8100
rect 2990 8195 3010 8215
rect 2990 8080 3010 8100
rect -3410 7900 -3390 7920
rect -3340 7900 -3320 7920
rect -2690 7900 -2670 7920
rect -2040 7900 -2020 7920
rect -1390 7900 -1370 7920
rect -740 7900 -720 7920
rect -30 6500 -10 6520
rect -125 5310 -105 5330
rect -125 5170 -105 5190
rect -125 2700 -105 2720
rect -85 2560 -65 2580
rect -55 1385 -35 1405
rect -3460 50 -3440 70
rect -3270 -30 -3250 -10
rect -3270 -160 -3250 -140
rect -2620 -30 -2600 -10
rect -2620 -160 -2600 -140
rect -1970 -30 -1950 -10
rect -1970 -160 -1950 -140
rect -1320 -30 -1300 -10
rect -1320 -160 -1300 -140
rect -670 -30 -650 -10
rect -670 -160 -650 -140
rect 515 -30 535 -10
rect 515 -160 535 -140
rect 1165 -30 1185 -10
rect 1165 -160 1185 -140
rect 1815 -30 1835 -10
rect 1815 -160 1835 -140
rect 2465 -30 2485 -10
rect 2465 -160 2485 -140
rect 3115 -30 3135 -10
rect 3115 -160 3135 -140
<< metal1 >>
rect -3530 -130 -3500 8225
rect -3460 7930 -3430 8225
rect -2520 8215 -2480 8225
rect -1870 8215 -1830 8225
rect -1220 8215 -1180 8225
rect -570 8215 -530 8225
rect 1030 8215 1070 8225
rect 1680 8215 1720 8225
rect 2330 8215 2370 8225
rect 2980 8215 3020 8225
rect -3165 8195 -2510 8215
rect -2490 8195 -1860 8215
rect -1840 8195 -1210 8215
rect -1190 8195 -560 8215
rect -540 8195 1040 8215
rect 1060 8195 1690 8215
rect 1710 8195 2340 8215
rect 2360 8195 2990 8215
rect 3010 8195 3280 8215
rect -3165 8185 3280 8195
rect -3460 7920 -3380 7930
rect -3460 7900 -3410 7920
rect -3390 7900 -3380 7920
rect -3460 7890 -3380 7900
rect -3350 7920 -3310 7930
rect -3350 7900 -3340 7920
rect -3320 7900 -3310 7920
rect -3350 7890 -3310 7900
rect -3165 7890 -3135 8185
rect -2950 8125 3280 8155
rect -2950 7890 -2920 8125
rect -2520 8100 -2480 8110
rect -2520 8080 -2510 8100
rect -2490 8080 -2480 8100
rect -2520 8070 -2480 8080
rect -2700 7920 -2660 7930
rect -2700 7900 -2690 7920
rect -2670 7900 -2660 7920
rect -2700 7890 -2660 7900
rect -2515 7890 -2485 8070
rect -2300 7890 -2270 8125
rect -1870 8100 -1830 8110
rect -1870 8080 -1860 8100
rect -1840 8080 -1830 8100
rect -1870 8070 -1830 8080
rect -2050 8020 -2010 8030
rect -2050 8000 -2040 8020
rect -2020 8000 -2010 8020
rect -2050 7990 -2010 8000
rect -2025 7930 -2010 7990
rect -2050 7920 -2010 7930
rect -2050 7900 -2040 7920
rect -2020 7900 -2010 7920
rect -2050 7890 -2010 7900
rect -1865 7890 -1835 8070
rect -1650 7890 -1620 8125
rect -1220 8100 -1180 8110
rect -1220 8080 -1210 8100
rect -1190 8080 -1180 8100
rect -1220 8070 -1180 8080
rect -1400 8060 -1360 8070
rect -1400 8040 -1390 8060
rect -1370 8040 -1360 8060
rect -1400 8030 -1360 8040
rect -1375 7930 -1360 8030
rect -1400 7920 -1360 7930
rect -1400 7900 -1390 7920
rect -1370 7900 -1360 7920
rect -1400 7890 -1360 7900
rect -1215 7890 -1185 8070
rect -1000 7890 -970 8125
rect -750 8100 -710 8110
rect -750 8080 -740 8100
rect -720 8080 -710 8100
rect -750 8070 -710 8080
rect -570 8100 -530 8110
rect -570 8080 -560 8100
rect -540 8080 -530 8100
rect -570 8070 -530 8080
rect -725 7930 -710 8070
rect -750 7920 -710 7930
rect -750 7900 -740 7920
rect -720 7900 -710 7920
rect -750 7890 -710 7900
rect -565 7890 -535 8070
rect -350 7890 -320 8125
rect 170 7890 200 8125
rect 820 7890 850 8125
rect 1030 8100 1070 8110
rect 1030 8080 1040 8100
rect 1060 8080 1070 8100
rect 1030 8070 1070 8080
rect 1035 7890 1065 8070
rect 1470 7890 1500 8125
rect 1680 8100 1720 8110
rect 1680 8080 1690 8100
rect 1710 8080 1720 8100
rect 1680 8070 1720 8080
rect 1685 7890 1715 8070
rect 2120 7890 2150 8125
rect 2330 8100 2370 8110
rect 2330 8080 2340 8100
rect 2360 8080 2370 8100
rect 2330 8070 2370 8080
rect 2335 7890 2365 8070
rect 2770 7890 2800 8125
rect 2980 8100 3020 8110
rect 2980 8080 2990 8100
rect 3010 8080 3020 8100
rect 2980 8070 3020 8080
rect 2985 7890 3015 8070
rect -3460 6615 -3430 7890
rect -3460 6575 -3400 6615
rect -3460 5300 -3430 6575
rect -40 6520 0 6530
rect -40 6500 -30 6520
rect -10 6500 0 6520
rect -40 6490 0 6500
rect -135 5330 -95 5340
rect -135 5310 -125 5330
rect -105 5315 -95 5330
rect -105 5310 -65 5315
rect -135 5300 -65 5310
rect -3460 5260 -3400 5300
rect -3460 3985 -3430 5260
rect -135 5190 -95 5200
rect -135 5170 -125 5190
rect -105 5170 -95 5190
rect -135 5160 -95 5170
rect -3460 3945 -3400 3985
rect -3460 2670 -3430 3945
rect -135 2730 -120 5160
rect -135 2720 -95 2730
rect -135 2700 -125 2720
rect -105 2700 -95 2720
rect -135 2690 -95 2700
rect -3460 2630 -3400 2670
rect -3460 1355 -3430 2630
rect -80 2590 -65 5300
rect -95 2580 -55 2590
rect -95 2560 -85 2580
rect -65 2560 -55 2580
rect -95 2550 -55 2560
rect -40 1415 -25 6490
rect -65 1405 -25 1415
rect -65 1385 -55 1405
rect -35 1385 -25 1405
rect -65 1375 -25 1385
rect -3460 1315 -3400 1355
rect -3460 80 -3430 1315
rect -3470 70 -3430 80
rect -3470 50 -3460 70
rect -3440 50 -3430 70
rect -3470 40 -3430 50
rect -3460 0 -3400 40
rect -3460 -70 -3430 0
rect -3285 -10 -3240 0
rect -3285 -30 -3270 -10
rect -3250 -30 -3240 -10
rect -3280 -40 -3240 -30
rect -3225 -70 -3195 0
rect -2795 -70 -2765 0
rect -2635 -10 -2590 0
rect -2635 -30 -2620 -10
rect -2600 -30 -2590 -10
rect -2630 -40 -2590 -30
rect -2575 -70 -2545 0
rect -2145 -70 -2115 0
rect -1985 -10 -1940 0
rect -1985 -30 -1970 -10
rect -1950 -30 -1940 -10
rect -1980 -40 -1940 -30
rect -1925 -70 -1895 0
rect -1495 -70 -1465 0
rect -1335 -10 -1290 0
rect -1335 -30 -1320 -10
rect -1300 -30 -1290 -10
rect -1330 -40 -1290 -30
rect -1275 -70 -1245 0
rect -845 -70 -815 0
rect -685 -10 -640 0
rect -685 -30 -670 -10
rect -650 -30 -640 -10
rect -680 -40 -640 -30
rect -625 -70 -595 0
rect -195 -70 -165 0
rect 15 -70 45 0
rect 445 -70 475 0
rect 505 -10 545 0
rect 505 -30 515 -10
rect 535 -30 545 -10
rect 505 -40 545 -30
rect 665 -70 695 0
rect 1095 -70 1125 0
rect 1155 -10 1195 0
rect 1155 -30 1165 -10
rect 1185 -30 1195 -10
rect 1155 -40 1195 -30
rect 1315 -70 1345 0
rect 1745 -70 1775 0
rect 1805 -10 1845 0
rect 1805 -30 1815 -10
rect 1835 -30 1845 -10
rect 1805 -40 1845 -30
rect 1965 -70 1995 0
rect 2395 -70 2425 0
rect 2455 -10 2495 0
rect 2455 -30 2465 -10
rect 2485 -30 2495 -10
rect 2455 -40 2495 -30
rect 2615 -70 2645 0
rect 3045 -70 3075 0
rect 3105 -10 3145 0
rect 3105 -30 3115 -10
rect 3135 -30 3145 -10
rect 3105 -40 3145 -30
rect 3250 -70 3280 7890
rect -3460 -100 3280 -70
rect -3530 -140 3280 -130
rect -3530 -160 -3270 -140
rect -3250 -160 -2620 -140
rect -2600 -160 -1970 -140
rect -1950 -160 -1320 -140
rect -1300 -160 -670 -140
rect -650 -160 515 -140
rect 535 -160 1165 -140
rect 1185 -160 1815 -140
rect 1835 -160 2465 -140
rect 2485 -160 3115 -140
rect 3135 -160 3280 -140
rect -3280 -170 -3240 -160
rect -2630 -170 -2590 -160
rect -1980 -170 -1940 -160
rect -1330 -170 -1290 -160
rect -680 -170 -640 -160
rect 505 -170 545 -160
rect 1155 -170 1195 -160
rect 1805 -170 1845 -160
rect 2455 -170 2495 -160
rect 3105 -170 3145 -160
use half_dac_for_mirroring  half_dac_for_mirroring_0
timestamp 1702420665
transform 1 0 650 0 1 1315
box -650 -1315 2600 6575
use half_dac_for_mirroring  half_dac_for_mirroring_1
timestamp 1702420665
transform -1 0 -800 0 -1 6575
box -650 -1315 2600 6575
<< labels >>
flabel locali -1960 8225 -1960 8225 1 FreeSans 160 0 0 0 X0
port 1 n
flabel locali -2000 8225 -2000 8225 1 FreeSans 160 0 0 0 X1
port 2 n
flabel locali -2040 8225 -2040 8225 1 FreeSans 160 0 0 0 X2
port 3 n
flabel locali -2080 8225 -2080 8225 1 FreeSans 160 0 0 0 X3
port 4 n
flabel locali -3450 8225 -3450 8225 1 FreeSans 160 0 0 0 Y0
port 5 n
flabel locali -3490 8225 -3490 8225 1 FreeSans 160 0 0 0 Y1
port 6 n
flabel locali -3530 8225 -3530 8225 1 FreeSans 160 0 0 0 Y2
port 7 n
flabel locali -3570 8225 -3570 8225 1 FreeSans 160 0 0 0 Y3
port 8 n
flabel metal1 3280 8140 3280 8140 3 FreeSans 160 0 0 0 I1
port 9 e
flabel metal1 3280 8200 3280 8200 3 FreeSans 160 0 0 0 I2
port 10 e
flabel metal1 3280 -145 3280 -145 3 FreeSans 160 0 0 0 VDD
port 11 e
flabel metal1 3280 -85 3280 -85 3 FreeSans 160 0 0 0 GND
port 12 e
<< end >>
