magic
tech sky130A
timestamp 1702744874
<< end >>
