magic
tech sky130A
timestamp 1702267426
<< nwell >>
rect 415 745 555 1225
<< nmos >>
rect 50 0 100 1200
rect 150 0 200 1200
rect 280 1140 380 1155
rect 280 1075 380 1090
rect 280 1010 380 1025
rect 280 815 380 830
rect 260 395 310 695
rect 260 0 310 300
<< pmos >>
rect 435 1140 535 1155
rect 435 1075 535 1090
rect 435 1010 535 1025
rect 435 815 535 830
<< ndiff >>
rect 0 0 50 1200
rect 100 0 150 1200
rect 200 695 250 1200
rect 280 1155 380 1205
rect 280 1090 380 1140
rect 280 1025 380 1075
rect 280 960 380 1010
rect 280 830 380 880
rect 280 765 380 815
rect 200 395 260 695
rect 310 395 360 695
rect 200 300 250 395
rect 200 0 260 300
rect 310 0 360 300
<< pdiff >>
rect 435 1155 535 1205
rect 435 1090 535 1140
rect 435 1025 535 1075
rect 435 960 535 1010
rect 435 830 535 880
rect 435 765 535 815
<< psubdiff >>
rect 280 915 380 930
rect 280 895 295 915
rect 365 895 380 915
rect 280 880 380 895
<< nsubdiff >>
rect 435 915 535 930
rect 435 895 450 915
rect 520 895 535 915
rect 435 880 535 895
<< psubdiffcont >>
rect 295 895 365 915
<< nsubdiffcont >>
rect 450 895 520 915
<< poly >>
rect 50 1200 100 1215
rect 150 1200 200 1215
rect 550 1165 590 1175
rect 550 1155 560 1165
rect 265 1140 280 1155
rect 380 1140 435 1155
rect 535 1145 560 1155
rect 580 1145 590 1165
rect 535 1140 590 1145
rect 550 1135 590 1140
rect 550 1100 590 1110
rect 550 1090 560 1100
rect 265 1075 280 1090
rect 380 1075 435 1090
rect 535 1080 560 1090
rect 580 1080 590 1100
rect 535 1075 590 1080
rect 550 1070 590 1075
rect 550 1035 590 1045
rect 550 1025 560 1035
rect 265 1010 280 1025
rect 380 1010 435 1025
rect 535 1015 560 1025
rect 580 1015 590 1035
rect 535 1010 590 1015
rect 550 1005 590 1010
rect 550 845 590 855
rect 550 830 560 845
rect 265 815 280 830
rect 380 815 435 830
rect 535 825 560 830
rect 580 825 590 845
rect 535 815 590 825
rect 260 740 310 750
rect 260 720 275 740
rect 295 720 310 740
rect 260 695 310 720
rect 260 380 310 395
rect 260 345 310 355
rect 260 325 275 345
rect 295 325 310 345
rect 260 300 310 325
rect 50 -15 100 0
rect 150 -15 200 0
rect 260 -15 310 0
<< polycont >>
rect 560 1145 580 1165
rect 560 1080 580 1100
rect 560 1015 580 1035
rect 560 825 580 845
rect 275 720 295 740
rect 275 325 295 345
<< locali >>
rect 0 1220 570 1240
rect 5 1185 45 1195
rect 5 15 15 1185
rect 35 15 45 1185
rect 285 1180 375 1200
rect 440 1180 530 1200
rect 245 1160 375 1180
rect 400 1160 530 1180
rect 550 1175 570 1220
rect 550 1165 590 1175
rect 245 1005 265 1160
rect 400 1070 420 1160
rect 550 1145 560 1165
rect 580 1145 590 1165
rect 550 1135 590 1145
rect 440 1125 530 1135
rect 440 1105 450 1125
rect 520 1105 530 1125
rect 440 1095 530 1105
rect 550 1100 590 1110
rect 550 1080 560 1100
rect 580 1080 590 1100
rect 550 1070 590 1080
rect 285 1060 375 1070
rect 285 1040 295 1060
rect 365 1040 375 1060
rect 400 1050 530 1070
rect 285 1030 375 1040
rect 440 1030 530 1050
rect 550 1035 590 1045
rect 550 1015 560 1035
rect 580 1015 590 1035
rect 550 1005 590 1015
rect 245 985 375 1005
rect 440 985 530 1005
rect 245 750 265 985
rect 285 965 570 985
rect 285 915 375 925
rect 285 895 295 915
rect 365 895 375 915
rect 285 865 375 895
rect 285 845 295 865
rect 365 845 375 865
rect 285 835 375 845
rect 440 915 530 925
rect 440 895 450 915
rect 520 895 530 915
rect 440 865 530 895
rect 440 845 450 865
rect 520 845 530 865
rect 440 835 530 845
rect 550 855 570 965
rect 550 845 590 855
rect 550 825 560 845
rect 580 825 590 845
rect 550 815 590 825
rect 285 790 375 810
rect 440 790 530 810
rect 285 770 530 790
rect 245 740 305 750
rect 245 730 275 740
rect 265 720 275 730
rect 295 720 305 740
rect 265 710 305 720
rect 315 680 355 690
rect 315 410 325 680
rect 345 410 355 680
rect 315 400 355 410
rect 375 355 395 770
rect 265 345 395 355
rect 265 325 275 345
rect 295 335 395 345
rect 295 325 305 335
rect 265 315 305 325
rect 5 5 45 15
rect 315 285 355 295
rect 315 15 325 285
rect 345 15 355 285
rect 315 5 355 15
<< viali >>
rect 15 15 35 1185
rect 450 1105 520 1125
rect 295 1040 365 1060
rect 295 895 365 915
rect 295 845 365 865
rect 450 895 520 915
rect 450 845 520 865
rect 325 410 345 680
rect 325 15 345 285
<< metal1 >>
rect 5 1185 45 1195
rect 5 15 15 1185
rect 35 15 45 1185
rect 285 1060 375 1240
rect 285 1040 295 1060
rect 365 1040 375 1060
rect 285 915 375 1040
rect 285 895 295 915
rect 365 895 375 915
rect 285 865 375 895
rect 285 845 295 865
rect 365 845 375 865
rect 285 835 375 845
rect 440 1125 530 1240
rect 440 1105 450 1125
rect 520 1105 530 1125
rect 440 915 530 1105
rect 440 895 450 915
rect 520 895 530 915
rect 440 865 530 895
rect 440 845 450 865
rect 520 845 530 865
rect 440 835 530 845
rect 315 680 355 690
rect 315 410 325 680
rect 345 410 355 680
rect 315 400 355 410
rect 5 5 45 15
rect 315 285 355 295
rect 315 15 325 285
rect 345 15 355 285
rect 315 5 355 15
<< end >>
