magic
tech sky130A
magscale 1 2
timestamp 1702679508
<< error_p >>
rect 3728 32860 3740 32862
rect 5028 32860 5040 32862
rect 6328 32860 6340 32862
rect 7628 32860 7640 32862
rect 8928 32860 8940 32862
rect 3750 32838 3752 32850
rect 5050 32838 5052 32850
rect 6350 32838 6352 32850
rect 7650 32838 7652 32850
rect 8950 32838 8952 32850
rect 10908 32140 10910 32152
rect 12208 32140 12210 32152
rect 13508 32140 13510 32152
rect 10920 32128 10932 32130
rect 12220 32128 12232 32130
rect 13520 32128 13532 32130
rect 3728 30230 3740 30232
rect 3750 30208 3752 30220
rect 9810 28630 9814 28650
rect 9776 28610 9780 28630
rect 3728 27600 3740 27602
rect 3750 27578 3752 27590
rect 3728 24970 3740 24972
rect 3750 24948 3752 24960
rect 3728 22340 3740 22342
rect 3750 22318 3752 22330
rect 3728 19710 3740 19712
rect 5028 19710 5040 19712
rect 6328 19710 6340 19712
rect 7628 19710 7640 19712
rect 8928 19710 8940 19712
rect 3750 19688 3752 19700
rect 5050 19688 5052 19700
rect 6350 19688 6352 19700
rect 7650 19688 7652 19700
rect 8950 19688 8952 19700
rect 10908 18990 10910 19002
rect 12208 18990 12210 19002
rect 13508 18990 13510 19002
rect 14808 18990 14810 19002
rect 10920 18978 10932 18980
rect 12220 18978 12232 18980
rect 13520 18978 13532 18980
rect 14820 18978 14832 18980
<< error_s >>
rect 16108 32140 16110 32152
rect 16120 32128 16132 32130
rect 16108 29510 16110 29522
rect 16120 29498 16132 29500
rect 16108 26880 16110 26892
rect 16120 26868 16132 26870
rect 16108 24250 16110 24262
rect 16120 24238 16132 24240
rect 16108 21620 16110 21632
rect 16120 21608 16132 21610
rect 16108 18990 16110 19002
rect 16120 18978 16132 18980
<< error_ps >>
rect 14808 32140 14810 32152
rect 14820 32128 14832 32130
<< locali >>
rect 2780 34680 2820 34820
rect 3460 34680 3500 34820
rect 2780 34660 2960 34680
rect 2780 34640 2900 34660
rect 2880 34620 2900 34640
rect 2940 34620 2960 34660
rect 2880 34600 2960 34620
rect 2920 34480 2960 34600
rect 3000 34640 3500 34680
rect 3000 34480 3040 34640
rect 3880 34600 3920 34820
rect 3080 34560 3920 34600
rect 3080 34480 3120 34560
rect 4140 34520 4180 34820
rect 4670 34740 4710 34820
rect 5350 34740 5390 34820
rect 5770 34740 5810 34820
rect 5900 34780 6070 34820
rect 4670 34720 4750 34740
rect 4670 34680 4690 34720
rect 4730 34680 4750 34720
rect 4670 34660 4750 34680
rect 5350 34720 5430 34740
rect 5350 34680 5370 34720
rect 5410 34680 5430 34720
rect 5350 34660 5430 34680
rect 5770 34720 5850 34740
rect 5770 34680 5790 34720
rect 5830 34680 5850 34720
rect 5770 34660 5850 34680
rect 3160 34480 4180 34520
rect 5900 34480 5940 34780
rect 5980 34720 6060 34740
rect 5980 34680 6000 34720
rect 6040 34680 6060 34720
rect 5980 34660 6060 34680
rect 5980 34480 6020 34660
rect 6100 34640 6180 34660
rect 6100 34620 6120 34640
rect 6060 34600 6120 34620
rect 6160 34600 6180 34640
rect 6060 34580 6180 34600
rect 6220 34580 6300 34600
rect 6060 34480 6100 34580
rect 6220 34540 6240 34580
rect 6280 34540 6300 34580
rect 6220 34520 6300 34540
rect 6140 34480 6260 34520
rect 19520 29150 19600 29170
rect 19520 29130 19540 29150
rect 19510 29110 19540 29130
rect 19580 29110 19600 29150
rect 19510 29090 19600 29110
rect 19510 27130 19710 27170
rect 19550 25080 19630 25100
rect 19550 25040 19570 25080
rect 19610 25040 19630 25080
rect 19550 25020 19630 25040
rect 19550 24500 19590 25020
rect 19510 24460 19590 24500
rect 19550 23680 19590 24460
rect 18200 23640 19590 23680
rect 18200 23530 18240 23640
rect 19670 23600 19710 27130
rect 18380 23560 19980 23600
rect 18380 23530 18420 23560
<< viali >>
rect 2900 34620 2940 34660
rect 4690 34680 4730 34720
rect 5370 34680 5410 34720
rect 5790 34680 5830 34720
rect 6000 34680 6040 34720
rect 6120 34600 6160 34640
rect 6240 34540 6280 34580
rect 19540 29110 19580 29150
rect 19570 25040 19610 25080
<< metal1 >>
rect 2880 34660 2960 34680
rect 2880 34620 2900 34660
rect 2940 34620 3080 34660
rect 2880 34600 3080 34620
rect 3020 34480 3080 34600
rect 3160 34480 3220 34850
rect 4670 34720 4750 34740
rect 4670 34680 4690 34720
rect 4730 34680 4750 34720
rect 4670 34660 4750 34680
rect 5350 34720 5430 34740
rect 5350 34680 5370 34720
rect 5410 34680 5430 34720
rect 5350 34660 5430 34680
rect 5770 34720 5850 34740
rect 5770 34680 5790 34720
rect 5830 34690 5850 34720
rect 5980 34720 6060 34740
rect 5980 34690 6000 34720
rect 5830 34680 6000 34690
rect 6040 34680 6060 34720
rect 5770 34660 6060 34680
rect 4720 34550 4750 34660
rect 5400 34610 5430 34660
rect 6100 34640 6180 34660
rect 6100 34610 6120 34640
rect 5400 34600 6120 34610
rect 6160 34600 6180 34640
rect 5400 34580 6180 34600
rect 6220 34580 6300 34600
rect 6220 34550 6240 34580
rect 4720 34540 6240 34550
rect 6280 34540 6300 34580
rect 4720 34520 6300 34540
rect 16640 34400 17770 34460
rect 16640 34280 17380 34340
rect 17320 33980 17380 34280
rect 17710 33900 17770 34400
rect 19550 31870 19600 31900
rect 19570 29170 19600 31870
rect 19520 29150 19600 29170
rect 19520 29110 19540 29150
rect 19580 29110 19600 29150
rect 19520 29090 19600 29110
rect 19550 25080 19630 25100
rect 19550 25040 19570 25080
rect 19610 25040 19630 25080
rect 19550 25020 19630 25040
rect 16700 23530 18200 23830
rect 18260 23650 19790 23680
rect 18260 23530 18290 23650
rect 18320 23590 20010 23620
rect 18320 23530 18350 23590
rect 16640 17830 16700 17890
rect 18420 17770 18480 17830
rect 16640 17710 18480 17770
use 4_bit_binary_decoder  4_bit_binary_decoder_0
timestamp 1702624819
transform 1 0 2780 0 1 34820
box -73 -54 3780 971
use bias  bias_0 ~/dev/git/magic-dds/magic
timestamp 1697165931
transform 0 1 16780 1 0 19350
box -1560 -150 4220 3210
use current_difference_balanced  current_difference_balanced_0
timestamp 1702677849
transform -1 0 19410 0 1 31510
box -140 -870 2680 2500
use current_steering_dac  current_steering_dac_0
timestamp 1702595941
transform 1 0 10080 0 1 18030
box -7300 -580 6560 16450
use opamp_balanced  opamp_balanced_0
timestamp 1702677968
transform -1 0 19410 0 1 24570
box -140 -870 2770 6050
<< end >>
