magic
tech sky130A
timestamp 1702371118
<< locali >>
rect -65 6505 0 6515
rect -65 6485 -55 6505
rect -35 6495 0 6505
rect -35 6485 -25 6495
rect -65 6475 -25 6485
rect -175 5330 -120 5340
rect -175 5320 -150 5330
rect -160 5310 -150 5320
rect -130 5310 -120 5330
rect -160 5300 -120 5310
rect -160 5190 0 5200
rect -160 5170 -150 5190
rect -130 5180 0 5190
rect -130 5170 -120 5180
rect -160 5160 -120 5170
rect -175 4005 -135 4025
rect -155 3885 -135 4005
rect -155 3865 0 3885
rect -160 2720 -120 2730
rect -160 2710 -150 2720
rect -175 2700 -150 2710
rect -130 2700 -120 2720
rect -175 2690 -120 2700
rect -120 2580 -80 2590
rect -120 2560 -110 2580
rect -90 2570 -80 2580
rect -90 2560 0 2570
rect -120 2550 0 2560
rect -90 1405 -50 1415
rect -90 1395 -80 1405
rect -175 1385 -80 1395
rect -60 1385 -50 1405
rect -175 1375 -50 1385
<< viali >>
rect -55 6485 -35 6505
rect -150 5310 -130 5330
rect -150 5170 -130 5190
rect -150 2700 -130 2720
rect -110 2560 -90 2580
rect -80 1385 -60 1405
<< metal1 >>
rect -65 6505 -25 6515
rect -65 6485 -55 6505
rect -35 6485 -25 6505
rect -65 6475 -25 6485
rect -160 5330 -120 5340
rect -160 5310 -150 5330
rect -130 5315 -120 5330
rect -130 5310 -90 5315
rect -160 5300 -90 5310
rect -160 5190 -120 5200
rect -160 5170 -150 5190
rect -130 5170 -120 5190
rect -160 5160 -120 5170
rect -160 2730 -145 5160
rect -160 2720 -120 2730
rect -160 2700 -150 2720
rect -130 2700 -120 2720
rect -160 2690 -120 2700
rect -105 2590 -90 5300
rect -120 2580 -80 2590
rect -120 2560 -110 2580
rect -90 2560 -80 2580
rect -120 2550 -80 2560
rect -65 1415 -50 6475
rect -90 1405 -50 1415
rect -90 1385 -80 1405
rect -60 1385 -50 1405
rect -90 1375 -50 1385
use half_dac_for_mirroring  half_dac_for_mirroring_0
timestamp 1702367632
transform 1 0 650 0 1 1315
box -650 -1315 2600 6575
use half_dac_for_mirroring  half_dac_for_mirroring_1
timestamp 1702367632
transform -1 0 -825 0 -1 6575
box -650 -1315 2600 6575
<< end >>
