magic
tech sky130A
timestamp 1702704436
<< error_s >>
rect -3176 7415 -3170 7416
rect -2526 7415 -2520 7416
rect -1876 7415 -1870 7416
rect -1226 7415 -1220 7416
rect -576 7415 -570 7416
rect -3165 7404 -3164 7410
rect -2515 7404 -2514 7410
rect -1865 7404 -1864 7410
rect -1215 7404 -1214 7410
rect -565 7404 -564 7410
rect 414 7055 415 7061
rect 1064 7055 1065 7061
rect 1714 7055 1715 7061
rect 2364 7055 2365 7061
rect 3014 7055 3015 7061
rect 420 7049 426 7050
rect 1070 7049 1076 7050
rect 1720 7049 1726 7050
rect 2370 7049 2376 7050
rect 3020 7049 3026 7050
rect -3176 6100 -3170 6101
rect -3165 6089 -3164 6095
rect 3014 5740 3015 5746
rect 3020 5734 3026 5735
rect -135 5300 -133 5310
rect -152 5290 -150 5300
rect -3176 4785 -3170 4786
rect -3165 4774 -3164 4780
rect 3014 4425 3015 4431
rect 3020 4419 3026 4420
rect -3176 3470 -3170 3471
rect -3165 3459 -3164 3465
rect 3014 3110 3015 3116
rect 3020 3104 3026 3105
rect -3176 2155 -3170 2156
rect -3165 2144 -3164 2150
rect 3014 1795 3015 1801
rect 3020 1789 3026 1790
rect -3176 840 -3170 841
rect -2526 840 -2520 841
rect -1876 840 -1870 841
rect -1226 840 -1220 841
rect -576 840 -570 841
rect -3165 829 -3164 835
rect -2515 829 -2514 835
rect -1865 829 -1864 835
rect -1215 829 -1214 835
rect -565 829 -564 835
rect 414 480 415 486
rect 1064 480 1065 486
rect 1714 480 1715 486
rect 2364 480 2365 486
rect 3014 480 3015 486
rect 420 474 426 475
rect 1070 474 1076 475
rect 1720 474 1726 475
rect 2370 474 2376 475
rect 3020 474 3026 475
<< poly >>
rect -2950 -10 -2900 0
rect -2950 -30 -2935 -10
rect -2915 -30 -2900 -10
rect -2950 -40 -2900 -30
rect -2850 -10 -2800 0
rect -2850 -30 -2835 -10
rect -2815 -30 -2800 -10
rect -2850 -40 -2800 -30
rect -2300 -10 -2250 0
rect -2300 -30 -2285 -10
rect -2265 -30 -2250 -10
rect -2300 -40 -2250 -30
rect -2200 -10 -2150 0
rect -2200 -30 -2185 -10
rect -2165 -30 -2150 -10
rect -2200 -40 -2150 -30
rect -1650 -10 -1600 0
rect -1650 -30 -1635 -10
rect -1615 -30 -1600 -10
rect -1650 -40 -1600 -30
rect -1550 -10 -1500 0
rect -1550 -30 -1535 -10
rect -1515 -30 -1500 -10
rect -1550 -40 -1500 -30
rect -1000 -10 -950 0
rect -1000 -30 -985 -10
rect -965 -30 -950 -10
rect -1000 -40 -950 -30
rect -900 -10 -850 0
rect -900 -30 -885 -10
rect -865 -30 -850 -10
rect -900 -40 -850 -30
rect -350 -10 -300 0
rect -350 -30 -335 -10
rect -315 -30 -300 -10
rect -350 -40 -300 -30
rect -250 -10 -200 0
rect -250 -30 -235 -10
rect -215 -30 -200 -10
rect -250 -40 -200 -30
rect 50 -10 100 0
rect 50 -30 65 -10
rect 85 -30 100 -10
rect 50 -40 100 -30
rect 150 -10 200 0
rect 150 -30 165 -10
rect 185 -30 200 -10
rect 150 -40 200 -30
rect 700 -10 750 0
rect 700 -30 715 -10
rect 735 -30 750 -10
rect 700 -40 750 -30
rect 800 -10 850 0
rect 800 -30 815 -10
rect 835 -30 850 -10
rect 800 -40 850 -30
rect 1350 -10 1400 0
rect 1350 -30 1365 -10
rect 1385 -30 1400 -10
rect 1350 -40 1400 -30
rect 1450 -10 1500 0
rect 1450 -30 1465 -10
rect 1485 -30 1500 -10
rect 1450 -40 1500 -30
rect 2000 -10 2050 0
rect 2000 -30 2015 -10
rect 2035 -30 2050 -10
rect 2000 -40 2050 -30
rect 2100 -10 2150 0
rect 2100 -30 2115 -10
rect 2135 -30 2150 -10
rect 2100 -40 2150 -30
rect 2650 -10 2700 0
rect 2650 -30 2665 -10
rect 2685 -30 2700 -10
rect 2650 -40 2700 -30
rect 2750 -10 2800 0
rect 2750 -30 2765 -10
rect 2785 -30 2800 -10
rect 2750 -40 2800 -30
<< polycont >>
rect -2935 -30 -2915 -10
rect -2835 -30 -2815 -10
rect -2285 -30 -2265 -10
rect -2185 -30 -2165 -10
rect -1635 -30 -1615 -10
rect -1535 -30 -1515 -10
rect -985 -30 -965 -10
rect -885 -30 -865 -10
rect -335 -30 -315 -10
rect -235 -30 -215 -10
rect 65 -30 85 -10
rect 165 -30 185 -10
rect 715 -30 735 -10
rect 815 -30 835 -10
rect 1365 -30 1385 -10
rect 1465 -30 1485 -10
rect 2015 -30 2035 -10
rect 2115 -30 2135 -10
rect 2665 -30 2685 -10
rect 2765 -30 2785 -10
<< locali >>
rect -3580 1395 -3560 8225
rect -3540 2710 -3520 8225
rect -3500 4025 -3480 8225
rect -3460 5340 -3440 8225
rect -2520 8215 -2480 8225
rect -2520 8195 -2510 8215
rect -2490 8195 -2480 8215
rect -2520 8100 -2480 8195
rect -2520 8080 -2510 8100
rect -2490 8080 -2480 8100
rect -2520 8070 -2480 8080
rect -2090 7970 -2070 8225
rect -2050 8030 -2030 8225
rect -2010 8070 -1990 8225
rect -1970 8110 -1950 8225
rect -1870 8215 -1830 8225
rect -1870 8195 -1860 8215
rect -1840 8195 -1830 8215
rect -1970 8090 -1930 8110
rect -2010 8050 -1970 8070
rect -2050 8020 -2010 8030
rect -2050 8000 -2040 8020
rect -2020 8000 -2010 8020
rect -2050 7990 -2010 8000
rect -1990 8010 -1970 8050
rect -1950 8050 -1930 8090
rect -1870 8100 -1830 8195
rect -1220 8215 -1180 8225
rect -1220 8195 -1210 8215
rect -1190 8195 -1180 8215
rect -1870 8080 -1860 8100
rect -1840 8080 -1830 8100
rect -1870 8070 -1830 8080
rect -1560 8090 -1320 8110
rect -1560 8050 -1540 8090
rect -1400 8060 -1360 8070
rect -1400 8050 -1390 8060
rect -1950 8030 -1540 8050
rect -1520 8040 -1390 8050
rect -1370 8040 -1360 8060
rect -1520 8030 -1360 8040
rect -1340 8050 -1320 8090
rect -1220 8100 -1180 8195
rect -570 8215 -530 8225
rect -570 8195 -560 8215
rect -540 8195 -530 8215
rect -1220 8080 -1210 8100
rect -1190 8080 -1180 8100
rect -1220 8070 -1180 8080
rect -910 8100 -710 8110
rect -910 8090 -740 8100
rect -910 8050 -890 8090
rect -750 8080 -740 8090
rect -720 8080 -710 8100
rect -750 8070 -710 8080
rect -570 8100 -530 8195
rect -570 8080 -560 8100
rect -540 8080 -530 8100
rect -570 8070 -530 8080
rect 380 8215 420 8225
rect 380 8195 390 8215
rect 410 8195 420 8215
rect 380 8100 420 8195
rect 380 8080 390 8100
rect 410 8080 420 8100
rect 380 8070 420 8080
rect 1030 8215 1070 8225
rect 1030 8195 1040 8215
rect 1060 8195 1070 8215
rect 1030 8100 1070 8195
rect 1030 8080 1040 8100
rect 1060 8080 1070 8100
rect 1030 8070 1070 8080
rect 1680 8215 1720 8225
rect 1680 8195 1690 8215
rect 1710 8195 1720 8215
rect 1680 8100 1720 8195
rect 1680 8080 1690 8100
rect 1710 8080 1720 8100
rect 1680 8070 1720 8080
rect 2330 8215 2370 8225
rect 2330 8195 2340 8215
rect 2360 8195 2370 8215
rect 2330 8100 2370 8195
rect 2330 8080 2340 8100
rect 2360 8080 2370 8100
rect 2330 8070 2370 8080
rect 2980 8215 3020 8225
rect 2980 8195 2990 8215
rect 3010 8195 3020 8215
rect 2980 8100 3020 8195
rect 2980 8080 2990 8100
rect 3010 8080 3020 8100
rect 2980 8070 3020 8080
rect -1340 8030 -890 8050
rect -870 8030 140 8050
rect -1520 8010 -1500 8030
rect -870 8010 -850 8030
rect 120 8010 140 8030
rect -1990 7990 -1500 8010
rect -1480 7990 -850 8010
rect -830 7990 100 8010
rect 120 7990 710 8010
rect -1480 7970 -1460 7990
rect -830 7970 -810 7990
rect 80 7970 100 7990
rect 690 7970 710 7990
rect -2090 7950 -1460 7970
rect -1440 7950 -810 7970
rect -790 7950 60 7970
rect 80 7950 670 7970
rect 690 7950 1320 7970
rect -2090 7930 -2070 7950
rect -1440 7930 -1420 7950
rect -790 7930 -770 7950
rect 40 7930 60 7950
rect 650 7930 670 7950
rect 1300 7930 1320 7950
rect -3420 7920 -3380 7930
rect -3420 7900 -3410 7920
rect -3390 7900 -3380 7920
rect -3420 7890 -3380 7900
rect -3350 7920 -3310 7930
rect -3350 7900 -3340 7920
rect -3320 7900 -3310 7920
rect -3350 7890 -3310 7900
rect -2700 7920 -2070 7930
rect -2700 7900 -2690 7920
rect -2670 7910 -2070 7920
rect -2050 7920 -1420 7930
rect -2670 7900 -2660 7910
rect -2700 7890 -2660 7900
rect -2050 7900 -2040 7920
rect -2020 7910 -1420 7920
rect -1400 7920 -770 7930
rect -2020 7900 -2010 7910
rect -2050 7890 -2010 7900
rect -1400 7900 -1390 7920
rect -1370 7910 -770 7920
rect -750 7920 0 7930
rect -1370 7900 -1360 7910
rect -1400 7890 -1360 7900
rect -750 7900 -740 7920
rect -720 7910 0 7920
rect 40 7910 630 7930
rect 650 7910 1280 7930
rect 1300 7910 1930 7930
rect -720 7900 -710 7910
rect -750 7890 -710 7900
rect -3420 6655 -3400 7890
rect -20 7850 0 7910
rect 610 7890 630 7910
rect 1260 7890 1280 7910
rect 1910 7890 1930 7910
rect -130 7810 0 7830
rect -130 6655 -110 7810
rect -3420 6635 -3380 6655
rect -150 6635 -110 6655
rect -60 6505 0 6515
rect -60 6485 -50 6505
rect -30 6495 0 6505
rect -30 6485 -20 6495
rect -60 6475 -20 6485
rect -3460 5320 -3380 5340
rect -150 5330 -95 5340
rect -150 5320 -125 5330
rect -135 5310 -125 5320
rect -105 5310 -95 5330
rect -135 5300 -95 5310
rect -135 5190 0 5200
rect -135 5170 -125 5190
rect -105 5180 0 5190
rect -105 5170 -95 5180
rect -135 5160 -95 5170
rect -3500 4005 -3380 4025
rect -150 4005 -110 4025
rect -130 3885 -110 4005
rect -130 3865 0 3885
rect -135 2720 -95 2730
rect -135 2710 -125 2720
rect -3540 2690 -3380 2710
rect -150 2700 -125 2710
rect -105 2700 -95 2720
rect -150 2690 -95 2700
rect -95 2580 -55 2590
rect -95 2560 -85 2580
rect -65 2570 -55 2580
rect -65 2560 0 2570
rect -95 2550 0 2560
rect -65 1405 -25 1415
rect -65 1395 -55 1405
rect -3580 1375 -3380 1395
rect -150 1385 -55 1395
rect -35 1385 -25 1405
rect -150 1375 -25 1385
rect -130 1235 0 1255
rect -130 80 -110 1235
rect -3470 70 -3380 80
rect -3470 50 -3460 70
rect -3440 60 -3380 70
rect -150 60 -110 80
rect -3440 50 -3430 60
rect -3470 40 -3430 50
rect -3280 -10 -3240 0
rect -3280 -30 -3270 -10
rect -3250 -30 -3240 -10
rect -3280 -140 -3240 -30
rect -3280 -160 -3270 -140
rect -3250 -160 -3240 -140
rect -3280 -170 -3240 -160
rect -2945 -10 -2905 0
rect -2945 -30 -2935 -10
rect -2915 -30 -2905 -10
rect -2945 -260 -2905 -30
rect -2845 -10 -2805 0
rect -2845 -30 -2835 -10
rect -2815 -30 -2805 -10
rect -2845 -200 -2805 -30
rect -2630 -10 -2590 0
rect -2630 -30 -2620 -10
rect -2600 -30 -2590 -10
rect -2630 -140 -2590 -30
rect -2630 -160 -2620 -140
rect -2600 -160 -2590 -140
rect -2630 -170 -2590 -160
rect -2295 -10 -2255 0
rect -2295 -30 -2285 -10
rect -2265 -30 -2255 -10
rect -2845 -220 -2835 -200
rect -2815 -220 -2805 -200
rect -2845 -230 -2805 -220
rect -2945 -280 -2935 -260
rect -2915 -280 -2905 -260
rect -2945 -290 -2905 -280
rect -2295 -260 -2255 -30
rect -2195 -10 -2155 0
rect -2195 -30 -2185 -10
rect -2165 -30 -2155 -10
rect -2195 -200 -2155 -30
rect -1980 -10 -1940 0
rect -1980 -30 -1970 -10
rect -1950 -30 -1940 -10
rect -1980 -140 -1940 -30
rect -1980 -160 -1970 -140
rect -1950 -160 -1940 -140
rect -1980 -170 -1940 -160
rect -1645 -10 -1605 0
rect -1645 -30 -1635 -10
rect -1615 -30 -1605 -10
rect -2195 -220 -2185 -200
rect -2165 -220 -2155 -200
rect -2195 -230 -2155 -220
rect -2295 -280 -2285 -260
rect -2265 -280 -2255 -260
rect -2295 -290 -2255 -280
rect -1645 -260 -1605 -30
rect -1545 -10 -1505 0
rect -1545 -30 -1535 -10
rect -1515 -30 -1505 -10
rect -1545 -200 -1505 -30
rect -1330 -10 -1290 0
rect -1330 -30 -1320 -10
rect -1300 -30 -1290 -10
rect -1330 -140 -1290 -30
rect -1330 -160 -1320 -140
rect -1300 -160 -1290 -140
rect -1330 -170 -1290 -160
rect -995 -10 -955 0
rect -995 -30 -985 -10
rect -965 -30 -955 -10
rect -1545 -220 -1535 -200
rect -1515 -220 -1505 -200
rect -1545 -230 -1505 -220
rect -1645 -280 -1635 -260
rect -1615 -280 -1605 -260
rect -1645 -290 -1605 -280
rect -995 -260 -955 -30
rect -895 -10 -855 0
rect -895 -30 -885 -10
rect -865 -30 -855 -10
rect -895 -200 -855 -30
rect -680 -10 -640 0
rect -680 -30 -670 -10
rect -650 -30 -640 -10
rect -680 -140 -640 -30
rect -680 -160 -670 -140
rect -650 -160 -640 -140
rect -680 -170 -640 -160
rect -345 -10 -305 0
rect -345 -30 -335 -10
rect -315 -30 -305 -10
rect -895 -220 -885 -200
rect -865 -220 -855 -200
rect -895 -230 -855 -220
rect -995 -280 -985 -260
rect -965 -280 -955 -260
rect -995 -290 -955 -280
rect -345 -260 -305 -30
rect -245 -10 -205 0
rect -245 -30 -235 -10
rect -215 -30 -205 -10
rect -245 -200 -205 -30
rect -245 -220 -235 -200
rect -215 -220 -205 -200
rect -245 -230 -205 -220
rect 55 -10 95 0
rect 55 -30 65 -10
rect 85 -30 95 -10
rect 55 -200 95 -30
rect 55 -220 65 -200
rect 85 -220 95 -200
rect 55 -230 95 -220
rect 155 -10 195 0
rect 155 -30 165 -10
rect 185 -30 195 -10
rect -345 -280 -335 -260
rect -315 -280 -305 -260
rect -345 -290 -305 -280
rect 155 -260 195 -30
rect 505 -10 545 0
rect 505 -30 515 -10
rect 535 -30 545 -10
rect 505 -140 545 -30
rect 505 -160 515 -140
rect 535 -160 545 -140
rect 505 -170 545 -160
rect 705 -10 745 0
rect 705 -30 715 -10
rect 735 -30 745 -10
rect 705 -200 745 -30
rect 705 -220 715 -200
rect 735 -220 745 -200
rect 705 -230 745 -220
rect 805 -10 845 0
rect 805 -30 815 -10
rect 835 -30 845 -10
rect 155 -280 165 -260
rect 185 -280 195 -260
rect 155 -290 195 -280
rect 805 -260 845 -30
rect 1155 -10 1195 0
rect 1155 -30 1165 -10
rect 1185 -30 1195 -10
rect 1155 -140 1195 -30
rect 1155 -160 1165 -140
rect 1185 -160 1195 -140
rect 1155 -170 1195 -160
rect 1355 -10 1395 0
rect 1355 -30 1365 -10
rect 1385 -30 1395 -10
rect 1355 -200 1395 -30
rect 1355 -220 1365 -200
rect 1385 -220 1395 -200
rect 1355 -230 1395 -220
rect 1455 -10 1495 0
rect 1455 -30 1465 -10
rect 1485 -30 1495 -10
rect 805 -280 815 -260
rect 835 -280 845 -260
rect 805 -290 845 -280
rect 1455 -260 1495 -30
rect 1805 -10 1845 0
rect 1805 -30 1815 -10
rect 1835 -30 1845 -10
rect 1805 -140 1845 -30
rect 1805 -160 1815 -140
rect 1835 -160 1845 -140
rect 1805 -170 1845 -160
rect 2005 -10 2045 0
rect 2005 -30 2015 -10
rect 2035 -30 2045 -10
rect 2005 -200 2045 -30
rect 2005 -220 2015 -200
rect 2035 -220 2045 -200
rect 2005 -230 2045 -220
rect 2105 -10 2145 0
rect 2105 -30 2115 -10
rect 2135 -30 2145 -10
rect 1455 -280 1465 -260
rect 1485 -280 1495 -260
rect 1455 -290 1495 -280
rect 2105 -260 2145 -30
rect 2455 -10 2495 0
rect 2455 -30 2465 -10
rect 2485 -30 2495 -10
rect 2455 -140 2495 -30
rect 2455 -160 2465 -140
rect 2485 -160 2495 -140
rect 2455 -170 2495 -160
rect 2655 -10 2695 0
rect 2655 -30 2665 -10
rect 2685 -30 2695 -10
rect 2655 -200 2695 -30
rect 2655 -220 2665 -200
rect 2685 -220 2695 -200
rect 2655 -230 2695 -220
rect 2755 -10 2795 0
rect 2755 -30 2765 -10
rect 2785 -30 2795 -10
rect 2105 -280 2115 -260
rect 2135 -280 2145 -260
rect 2105 -290 2145 -280
rect 2755 -260 2795 -30
rect 3105 -10 3145 0
rect 3105 -30 3115 -10
rect 3135 -30 3145 -10
rect 3105 -140 3145 -30
rect 3105 -160 3115 -140
rect 3135 -160 3145 -140
rect 3105 -170 3145 -160
rect 2755 -280 2765 -260
rect 2785 -280 2795 -260
rect 2755 -290 2795 -280
<< viali >>
rect -2510 8195 -2490 8215
rect -2510 8080 -2490 8100
rect -1860 8195 -1840 8215
rect -2040 8000 -2020 8020
rect -1210 8195 -1190 8215
rect -1860 8080 -1840 8100
rect -1390 8040 -1370 8060
rect -560 8195 -540 8215
rect -1210 8080 -1190 8100
rect -740 8080 -720 8100
rect -560 8080 -540 8100
rect 390 8195 410 8215
rect 390 8080 410 8100
rect 1040 8195 1060 8215
rect 1040 8080 1060 8100
rect 1690 8195 1710 8215
rect 1690 8080 1710 8100
rect 2340 8195 2360 8215
rect 2340 8080 2360 8100
rect 2990 8195 3010 8215
rect 2990 8080 3010 8100
rect -3410 7900 -3390 7920
rect -3340 7900 -3320 7920
rect -2690 7900 -2670 7920
rect -2040 7900 -2020 7920
rect -1390 7900 -1370 7920
rect -740 7900 -720 7920
rect -50 6485 -30 6505
rect -125 5310 -105 5330
rect -125 5170 -105 5190
rect -125 2700 -105 2720
rect -85 2560 -65 2580
rect -55 1385 -35 1405
rect -3460 50 -3440 70
rect -3270 -30 -3250 -10
rect -3270 -160 -3250 -140
rect -2620 -30 -2600 -10
rect -2620 -160 -2600 -140
rect -2835 -220 -2815 -200
rect -2935 -280 -2915 -260
rect -1970 -30 -1950 -10
rect -1970 -160 -1950 -140
rect -2185 -220 -2165 -200
rect -2285 -280 -2265 -260
rect -1320 -30 -1300 -10
rect -1320 -160 -1300 -140
rect -1535 -220 -1515 -200
rect -1635 -280 -1615 -260
rect -670 -30 -650 -10
rect -670 -160 -650 -140
rect -885 -220 -865 -200
rect -985 -280 -965 -260
rect -235 -220 -215 -200
rect 65 -220 85 -200
rect -335 -280 -315 -260
rect 515 -30 535 -10
rect 515 -160 535 -140
rect 715 -220 735 -200
rect 165 -280 185 -260
rect 1165 -30 1185 -10
rect 1165 -160 1185 -140
rect 1365 -220 1385 -200
rect 815 -280 835 -260
rect 1815 -30 1835 -10
rect 1815 -160 1835 -140
rect 2015 -220 2035 -200
rect 1465 -280 1485 -260
rect 2465 -30 2485 -10
rect 2465 -160 2485 -140
rect 2665 -220 2685 -200
rect 2115 -280 2135 -260
rect 3115 -30 3135 -10
rect 3115 -160 3135 -140
rect 2765 -280 2785 -260
<< metal1 >>
rect -3650 -260 -3620 8225
rect -3590 -200 -3560 8225
rect -3530 -130 -3500 8225
rect -3460 7930 -3430 8225
rect -2520 8215 -2480 8225
rect -1870 8215 -1830 8225
rect -1220 8215 -1180 8225
rect -570 8215 -530 8225
rect 380 8215 420 8225
rect 1030 8215 1070 8225
rect 1680 8215 1720 8225
rect 2330 8215 2370 8225
rect 2980 8215 3020 8225
rect -3165 8195 -2510 8215
rect -2490 8195 -1860 8215
rect -1840 8195 -1210 8215
rect -1190 8195 -560 8215
rect -540 8195 390 8215
rect 410 8195 1040 8215
rect 1060 8195 1690 8215
rect 1710 8195 2340 8215
rect 2360 8195 2990 8215
rect 3010 8195 3280 8215
rect -3165 8185 3280 8195
rect -3460 7920 -3310 7930
rect -3460 7900 -3410 7920
rect -3390 7900 -3340 7920
rect -3320 7900 -3310 7920
rect -3460 7890 -3310 7900
rect -3165 7890 -3135 8185
rect -2950 8125 3280 8155
rect -2950 7890 -2920 8125
rect -2520 8100 -2480 8110
rect -2520 8080 -2510 8100
rect -2490 8080 -2480 8100
rect -2520 8070 -2480 8080
rect -2700 7920 -2660 7930
rect -2700 7900 -2690 7920
rect -2670 7900 -2660 7920
rect -2700 7890 -2660 7900
rect -2515 7890 -2485 8070
rect -2300 7890 -2270 8125
rect -1870 8100 -1830 8110
rect -1870 8080 -1860 8100
rect -1840 8080 -1830 8100
rect -1870 8070 -1830 8080
rect -2050 8020 -2010 8030
rect -2050 8000 -2040 8020
rect -2020 8000 -2010 8020
rect -2050 7990 -2010 8000
rect -2025 7930 -2010 7990
rect -2050 7920 -2010 7930
rect -2050 7900 -2040 7920
rect -2020 7900 -2010 7920
rect -2050 7890 -2010 7900
rect -1865 7890 -1835 8070
rect -1650 7890 -1620 8125
rect -1220 8100 -1180 8110
rect -1220 8080 -1210 8100
rect -1190 8080 -1180 8100
rect -1220 8070 -1180 8080
rect -1400 8060 -1360 8070
rect -1400 8040 -1390 8060
rect -1370 8040 -1360 8060
rect -1400 8030 -1360 8040
rect -1375 7930 -1360 8030
rect -1400 7920 -1360 7930
rect -1400 7900 -1390 7920
rect -1370 7900 -1360 7920
rect -1400 7890 -1360 7900
rect -1215 7890 -1185 8070
rect -1000 7890 -970 8125
rect -750 8100 -710 8110
rect -750 8080 -740 8100
rect -720 8080 -710 8100
rect -750 8070 -710 8080
rect -570 8100 -530 8110
rect -570 8080 -560 8100
rect -540 8080 -530 8100
rect -570 8070 -530 8080
rect -725 7930 -710 8070
rect -750 7920 -710 7930
rect -750 7900 -740 7920
rect -720 7900 -710 7920
rect -750 7890 -710 7900
rect -565 7890 -535 8070
rect -350 7890 -320 8125
rect 170 7890 200 8125
rect 380 8100 420 8110
rect 380 8080 390 8100
rect 410 8080 420 8100
rect 380 8070 420 8080
rect 385 7890 415 8070
rect 820 7890 850 8125
rect 1030 8100 1070 8110
rect 1030 8080 1040 8100
rect 1060 8080 1070 8100
rect 1030 8070 1070 8080
rect 1035 7890 1065 8070
rect 1470 7890 1500 8125
rect 1680 8100 1720 8110
rect 1680 8080 1690 8100
rect 1710 8080 1720 8100
rect 1680 8070 1720 8080
rect 1685 7890 1715 8070
rect 2120 7890 2150 8125
rect 2330 8100 2370 8110
rect 2330 8080 2340 8100
rect 2360 8080 2370 8100
rect 2330 8070 2370 8080
rect 2335 7890 2365 8070
rect 2770 7890 2800 8125
rect 2980 8100 3020 8110
rect 2980 8080 2990 8100
rect 3010 8080 3020 8100
rect 2980 8070 3020 8080
rect 2985 7890 3015 8070
rect -3460 6615 -3430 7890
rect -3460 6575 -3400 6615
rect -3460 5300 -3430 6575
rect -60 6505 -20 6515
rect -60 6485 -50 6505
rect -30 6485 -20 6505
rect -60 6475 -20 6485
rect -135 5330 -95 5340
rect -135 5310 -125 5330
rect -105 5315 -95 5330
rect -105 5310 -65 5315
rect -135 5300 -65 5310
rect -3460 5260 -3400 5300
rect -3460 3985 -3430 5260
rect -135 5190 -95 5200
rect -135 5170 -125 5190
rect -105 5170 -95 5190
rect -135 5160 -95 5170
rect -3460 3945 -3400 3985
rect -3460 2670 -3430 3945
rect -135 2730 -120 5160
rect -135 2720 -95 2730
rect -135 2700 -125 2720
rect -105 2700 -95 2720
rect -135 2690 -95 2700
rect -3460 2630 -3400 2670
rect -3460 1355 -3430 2630
rect -80 2590 -65 5300
rect -95 2580 -55 2590
rect -95 2560 -85 2580
rect -65 2560 -55 2580
rect -95 2550 -55 2560
rect -40 1415 -25 6475
rect -65 1405 -25 1415
rect -65 1385 -55 1405
rect -35 1385 -25 1405
rect -65 1375 -25 1385
rect -3460 1315 -3400 1355
rect -3460 80 -3430 1315
rect -3470 70 -3430 80
rect -3470 50 -3460 70
rect -3440 50 -3430 70
rect -3470 40 -3430 50
rect -3460 0 -3400 40
rect -3460 -70 -3430 0
rect -3285 -10 -3240 0
rect -3285 -30 -3270 -10
rect -3250 -30 -3240 -10
rect -3280 -40 -3240 -30
rect -3225 -70 -3195 0
rect -2795 -70 -2765 0
rect -2635 -10 -2590 0
rect -2635 -30 -2620 -10
rect -2600 -30 -2590 -10
rect -2630 -40 -2590 -30
rect -2575 -70 -2545 0
rect -2145 -70 -2115 0
rect -1985 -10 -1940 0
rect -1985 -30 -1970 -10
rect -1950 -30 -1940 -10
rect -1980 -40 -1940 -30
rect -1925 -70 -1895 0
rect -1495 -70 -1465 0
rect -1335 -10 -1290 0
rect -1335 -30 -1320 -10
rect -1300 -30 -1290 -10
rect -1330 -40 -1290 -30
rect -1275 -70 -1245 0
rect -845 -70 -815 0
rect -685 -10 -640 0
rect -685 -30 -670 -10
rect -650 -30 -640 -10
rect -680 -40 -640 -30
rect -625 -70 -595 0
rect -195 -70 -165 0
rect 15 -70 45 0
rect 445 -70 475 0
rect 505 -10 545 0
rect 505 -30 515 -10
rect 535 -30 545 -10
rect 505 -40 545 -30
rect 665 -70 695 0
rect 1095 -70 1125 0
rect 1155 -10 1195 0
rect 1155 -30 1165 -10
rect 1185 -30 1195 -10
rect 1155 -40 1195 -30
rect 1315 -70 1345 0
rect 1745 -70 1775 0
rect 1805 -10 1845 0
rect 1805 -30 1815 -10
rect 1835 -30 1845 -10
rect 1805 -40 1845 -30
rect 1965 -70 1995 0
rect 2395 -70 2425 0
rect 2455 -10 2495 0
rect 2455 -30 2465 -10
rect 2485 -30 2495 -10
rect 2455 -40 2495 -30
rect 2615 -70 2645 0
rect 3045 -70 3075 0
rect 3105 -10 3145 0
rect 3105 -30 3115 -10
rect 3135 -30 3145 -10
rect 3105 -40 3145 -30
rect 3160 -70 3175 0
rect 3250 -70 3280 7890
rect -3460 -100 3280 -70
rect -3530 -140 3280 -130
rect -3530 -160 -3270 -140
rect -3250 -160 -2620 -140
rect -2600 -160 -1970 -140
rect -1950 -160 -1320 -140
rect -1300 -160 -670 -140
rect -650 -160 515 -140
rect 535 -160 1165 -140
rect 1185 -160 1815 -140
rect 1835 -160 2465 -140
rect 2485 -160 3115 -140
rect 3135 -160 3280 -140
rect -3280 -170 -3240 -160
rect -2630 -170 -2590 -160
rect -1980 -170 -1940 -160
rect -1330 -170 -1290 -160
rect -680 -170 -640 -160
rect 505 -170 545 -160
rect 1155 -170 1195 -160
rect 1805 -170 1845 -160
rect 2455 -170 2495 -160
rect 3105 -170 3145 -160
rect -2845 -200 -2805 -190
rect -2195 -200 -2155 -190
rect -1545 -200 -1505 -190
rect -895 -200 -855 -190
rect -245 -200 -205 -190
rect 55 -200 95 -190
rect 705 -200 745 -190
rect 1355 -200 1395 -190
rect 2005 -200 2045 -190
rect 2655 -200 2695 -190
rect -3590 -220 -2835 -200
rect -2815 -220 -2185 -200
rect -2165 -220 -1535 -200
rect -1515 -220 -885 -200
rect -865 -220 -235 -200
rect -215 -220 65 -200
rect 85 -220 715 -200
rect 735 -220 1365 -200
rect 1385 -220 2015 -200
rect 2035 -220 2665 -200
rect 2685 -220 3280 -200
rect -3590 -230 3280 -220
rect -2945 -260 -2905 -250
rect -2295 -260 -2255 -250
rect -1645 -260 -1605 -250
rect -995 -260 -955 -250
rect -345 -260 -305 -250
rect 155 -260 195 -250
rect 805 -260 845 -250
rect 1455 -260 1495 -250
rect 2105 -260 2145 -250
rect 2755 -260 2795 -250
rect -3650 -280 -2935 -260
rect -2915 -280 -2285 -260
rect -2265 -280 -1635 -260
rect -1615 -280 -985 -260
rect -965 -280 -335 -260
rect -315 -280 165 -260
rect 185 -280 815 -260
rect 835 -280 1465 -260
rect 1485 -280 2115 -260
rect 2135 -280 2765 -260
rect 2785 -280 3280 -260
rect -3650 -290 3280 -280
use half_dac_for_mirroring  half_dac_for_mirroring_0
timestamp 1702704436
transform 1 0 650 0 1 1315
box -698 -1315 2600 6575
use half_dac_for_mirroring  half_dac_for_mirroring_1
timestamp 1702704436
transform -1 0 -800 0 -1 6575
box -698 -1315 2600 6575
<< labels >>
flabel locali -1960 8225 -1960 8225 1 FreeSans 160 0 0 0 X0
port 1 n
flabel locali -2000 8225 -2000 8225 1 FreeSans 160 0 0 0 X1
port 2 n
flabel locali -2040 8225 -2040 8225 1 FreeSans 160 0 0 0 X2
port 3 n
flabel locali -2080 8225 -2080 8225 1 FreeSans 160 0 0 0 X3
port 4 n
flabel locali -3450 8225 -3450 8225 1 FreeSans 160 0 0 0 Y0
port 5 n
flabel locali -3490 8225 -3490 8225 1 FreeSans 160 0 0 0 Y1
port 6 n
flabel locali -3530 8225 -3530 8225 1 FreeSans 160 0 0 0 Y2
port 7 n
flabel locali -3570 8225 -3570 8225 1 FreeSans 160 0 0 0 Y3
port 8 n
flabel metal1 3280 8140 3280 8140 3 FreeSans 160 0 0 0 I1
port 9 e
flabel metal1 3280 8200 3280 8200 3 FreeSans 160 0 0 0 I2
port 10 e
flabel metal1 3280 -145 3280 -145 3 FreeSans 160 0 0 0 VDD
port 11 e
flabel metal1 3280 -85 3280 -85 3 FreeSans 160 0 0 0 GND
port 12 e
flabel metal1 3280 -215 3280 -215 3 FreeSans 240 0 0 0 Vbn
port 13 e
flabel metal1 3280 -275 3280 -275 3 FreeSans 240 0 0 0 Vcn
port 14 e
<< end >>
