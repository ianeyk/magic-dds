magic
tech sky130A
magscale 1 2
timestamp 1702789236
<< nwell >>
rect 20690 31640 20950 34120
<< xpolycontact >>
rect 16780 33480 16920 33920
rect 16780 30740 16920 31180
rect 17170 33480 17310 33920
rect 17170 30740 17310 31180
rect 17560 33480 17700 33920
rect 17560 30740 17700 31180
rect 17950 33480 18090 33920
rect 17950 30740 18090 31180
rect 18340 33480 18480 33920
rect 18340 30740 18480 31180
rect 18730 33480 18870 33920
rect 18730 30740 18870 31180
<< xpolyres >>
rect 16780 31180 16920 33480
rect 17170 31180 17310 33480
rect 17560 31180 17700 33480
rect 17950 31180 18090 33480
rect 18340 31180 18480 33480
rect 18730 31180 18870 33480
<< locali >>
rect 2780 34680 2820 34820
rect 3460 34680 3500 34820
rect 2780 34660 2960 34680
rect 2780 34640 2900 34660
rect 2880 34620 2900 34640
rect 2940 34620 2960 34660
rect 2880 34600 2960 34620
rect 2920 34480 2960 34600
rect 3000 34640 3500 34680
rect 3000 34480 3040 34640
rect 3880 34600 3920 34820
rect 3080 34560 3920 34600
rect 3080 34480 3120 34560
rect 4140 34520 4180 34820
rect 4670 34740 4710 34820
rect 5350 34740 5390 34820
rect 5770 34740 5810 34820
rect 5900 34780 6070 34820
rect 4670 34720 4750 34740
rect 4670 34680 4690 34720
rect 4730 34680 4750 34720
rect 4670 34660 4750 34680
rect 5350 34720 5430 34740
rect 5350 34680 5370 34720
rect 5410 34680 5430 34720
rect 5350 34660 5430 34680
rect 5770 34720 5850 34740
rect 5770 34680 5790 34720
rect 5830 34680 5850 34720
rect 5770 34660 5850 34680
rect 3160 34480 4180 34520
rect 5900 34480 5940 34780
rect 5980 34720 6060 34740
rect 5980 34680 6000 34720
rect 6040 34680 6060 34720
rect 5980 34660 6060 34680
rect 5980 34480 6020 34660
rect 6100 34640 6180 34660
rect 6100 34620 6120 34640
rect 6060 34600 6120 34620
rect 6160 34600 6180 34640
rect 6060 34580 6180 34600
rect 6220 34580 6300 34600
rect 6060 34480 6100 34580
rect 6220 34540 6240 34580
rect 6280 34540 6300 34580
rect 6220 34520 6300 34540
rect 6140 34480 6260 34520
rect 17170 34460 17250 34480
rect 17170 34420 17190 34460
rect 17230 34420 17250 34460
rect 16780 34320 16860 34340
rect 16780 34280 16800 34320
rect 16840 34280 16860 34320
rect 16780 33920 16860 34280
rect 17170 33920 17250 34420
rect 18010 34000 18810 34080
rect 18010 33920 18090 34000
rect 18730 33920 18810 34000
rect 17620 33400 17700 33480
rect 18340 33400 18420 33480
rect 17620 33320 18420 33400
rect 20480 31840 20560 34070
rect 20470 31820 20570 31840
rect 20470 31760 20490 31820
rect 20550 31760 20570 31820
rect 20470 31740 20570 31760
rect 16840 31270 17640 31340
rect 16840 31180 16920 31270
rect 17560 31180 17640 31270
rect 18400 31320 20140 31340
rect 18400 31280 19760 31320
rect 19800 31280 20140 31320
rect 18400 31260 20140 31280
rect 18400 31180 18480 31260
rect 18870 30840 20040 30860
rect 18870 30800 19980 30840
rect 20020 30800 20040 30840
rect 18870 30780 20040 30800
rect 20480 30780 20560 31740
rect 20840 30800 20880 30840
rect 20820 30740 20860 30780
rect 17230 30650 17310 30740
rect 17950 30650 18030 30740
rect 19870 30720 23520 30740
rect 19870 30680 19890 30720
rect 19930 30700 23520 30720
rect 19930 30680 19950 30700
rect 19870 30660 19950 30680
rect 17230 30580 18030 30650
rect 19510 30600 20350 30620
rect 19510 30580 19820 30600
rect 19800 30560 19820 30580
rect 19860 30580 20350 30600
rect 19860 30560 19880 30580
rect 19800 30540 19880 30560
rect 19570 30080 19650 30100
rect 19570 30060 19590 30080
rect 19510 30040 19590 30060
rect 19630 30040 19650 30080
rect 19510 30020 19650 30040
rect 19990 30080 20070 30100
rect 19990 30040 20010 30080
rect 20050 30060 20070 30080
rect 20050 30040 20130 30060
rect 19990 30020 20130 30040
rect 19500 29770 20360 29850
rect 19630 29190 19710 29210
rect 19630 29150 19650 29190
rect 19690 29150 19710 29190
rect 19630 29130 19710 29150
rect 19980 29150 20060 29170
rect 19510 29090 19670 29130
rect 19980 29110 20000 29150
rect 20040 29130 20060 29150
rect 20040 29110 20130 29130
rect 19980 29090 20130 29110
rect 20170 29090 20350 29130
rect 19510 28960 20350 28980
rect 19510 28940 19830 28960
rect 19810 28920 19830 28940
rect 19870 28940 20350 28960
rect 19870 28920 19890 28940
rect 19810 28900 19890 28920
rect 19500 27260 20360 27340
rect 19510 27130 20350 27170
rect 19670 25080 19710 27130
rect 19670 25060 19750 25080
rect 19670 25020 19690 25060
rect 19730 25020 19750 25060
rect 19670 25000 19750 25020
rect 19560 24940 19640 24960
rect 19560 24900 19580 24940
rect 19620 24900 19640 24940
rect 19560 24880 19640 24900
rect 19510 24460 20350 24500
rect 19550 23680 19590 24460
rect 18200 23640 19590 23680
rect 19670 23830 19770 23850
rect 19670 23790 19710 23830
rect 19750 23790 19770 23830
rect 19670 23770 19770 23790
rect 18200 23530 18240 23640
rect 19670 23600 19710 23770
rect 18380 23560 19710 23600
rect 19920 23740 20420 23760
rect 19920 23700 20360 23740
rect 20400 23700 20420 23740
rect 19920 23680 20420 23700
rect 18380 23530 18420 23560
rect 19920 23520 20000 23680
rect 20130 23590 21770 23600
rect 19890 23440 20000 23520
rect 20090 23570 21770 23590
rect 20090 23530 20110 23570
rect 20150 23560 21770 23570
rect 20150 23530 20170 23560
rect 21730 23530 21770 23560
rect 20090 23510 20170 23530
rect 18350 17450 18390 17830
rect 21880 17450 21920 17830
<< viali >>
rect 2900 34620 2940 34660
rect 4690 34680 4730 34720
rect 5370 34680 5410 34720
rect 5790 34680 5830 34720
rect 6000 34680 6040 34720
rect 6120 34600 6160 34640
rect 6240 34540 6280 34580
rect 17190 34420 17230 34460
rect 16800 34280 16840 34320
rect 20290 34010 20330 34050
rect 20710 34010 20750 34050
rect 20840 31860 20880 31900
rect 20490 31760 20550 31820
rect 19760 31280 19800 31320
rect 19980 30800 20020 30840
rect 20420 30800 20460 30840
rect 19890 30680 19930 30720
rect 19820 30560 19860 30600
rect 19590 30040 19630 30080
rect 20010 30040 20050 30080
rect 19650 29150 19690 29190
rect 20000 29110 20040 29150
rect 19830 28920 19870 28960
rect 19690 25020 19730 25060
rect 19580 24900 19620 24940
rect 19710 23790 19750 23830
rect 20360 23700 20400 23740
rect 20110 23530 20150 23570
<< metal1 >>
rect 2880 34660 2960 34680
rect 2880 34620 2900 34660
rect 2940 34620 3080 34660
rect 2880 34600 3080 34620
rect 3020 34480 3080 34600
rect 3160 34480 3220 34850
rect 4670 34720 4750 34740
rect 4670 34680 4690 34720
rect 4730 34680 4750 34720
rect 4670 34660 4750 34680
rect 5350 34720 5430 34740
rect 5350 34680 5370 34720
rect 5410 34680 5430 34720
rect 5350 34660 5430 34680
rect 5770 34720 5850 34740
rect 5770 34680 5790 34720
rect 5830 34690 5850 34720
rect 5980 34720 6060 34740
rect 5980 34690 6000 34720
rect 5830 34680 6000 34690
rect 6040 34680 6060 34720
rect 5770 34660 6060 34680
rect 4720 34550 4750 34660
rect 5400 34610 5430 34660
rect 6100 34640 6180 34660
rect 6100 34610 6120 34640
rect 5400 34600 6120 34610
rect 6160 34600 6180 34640
rect 5400 34580 6180 34600
rect 6220 34580 6300 34600
rect 6220 34550 6240 34580
rect 4720 34540 6240 34550
rect 6280 34540 6300 34580
rect 4720 34520 6300 34540
rect 17170 34460 17250 34480
rect 16640 34420 17190 34460
rect 17230 34420 19710 34460
rect 16640 34400 19710 34420
rect 16640 34320 19600 34340
rect 16640 34280 16800 34320
rect 16840 34280 19600 34320
rect 16780 34260 16860 34280
rect 19570 30100 19600 34280
rect 19570 30080 19650 30100
rect 19570 30040 19590 30080
rect 19630 30040 19650 30080
rect 19570 30020 19650 30040
rect 19680 29210 19710 34400
rect 19630 29190 19710 29210
rect 19630 29150 19650 29190
rect 19690 29150 19710 29190
rect 19630 29130 19710 29150
rect 19740 31930 19770 34460
rect 19740 31920 19870 31930
rect 19740 31840 19780 31920
rect 19860 31840 19870 31920
rect 19740 31830 19870 31840
rect 19740 31340 19770 31830
rect 19740 31320 19820 31340
rect 19740 31280 19760 31320
rect 19800 31280 19820 31320
rect 19740 31260 19820 31280
rect 19740 29100 19770 31260
rect 19980 30860 20010 35750
rect 20260 34390 20360 34400
rect 20260 34310 20270 34390
rect 20350 34310 20360 34390
rect 20260 34300 20360 34310
rect 20680 34390 20780 34400
rect 20680 34310 20690 34390
rect 20770 34310 20780 34390
rect 20680 34300 20780 34310
rect 20270 34050 20350 34300
rect 20270 34010 20290 34050
rect 20330 34010 20350 34050
rect 20270 33990 20350 34010
rect 20690 34050 20770 34300
rect 20690 34010 20710 34050
rect 20750 34010 20770 34050
rect 20690 33990 20770 34010
rect 20810 31920 20910 31930
rect 20810 31840 20820 31920
rect 20900 31840 20910 31920
rect 20470 31830 20570 31840
rect 20810 31830 20910 31840
rect 20470 31750 20480 31830
rect 20560 31750 20570 31830
rect 20470 31740 20570 31750
rect 19960 30840 20040 30860
rect 19960 30800 19980 30840
rect 20020 30800 20040 30840
rect 19960 30780 20040 30800
rect 20400 30840 20480 30860
rect 20400 30800 20420 30840
rect 20460 30800 20480 30840
rect 20400 30780 20480 30800
rect 19870 30720 19950 30740
rect 19870 30680 19890 30720
rect 19930 30680 19950 30720
rect 19870 30660 19950 30680
rect 19690 29070 19770 29100
rect 19800 30600 19880 30620
rect 19800 30560 19820 30600
rect 19860 30560 19880 30600
rect 19800 30540 19880 30560
rect 19690 28810 19720 29070
rect 19800 29040 19830 30540
rect 19920 30220 19950 30660
rect 19870 30190 19950 30220
rect 19870 29930 19900 30190
rect 19980 30160 20010 30780
rect 20400 30750 20430 30780
rect 19930 30130 20010 30160
rect 20040 30720 20430 30750
rect 19930 29990 19960 30130
rect 20040 30100 20070 30720
rect 19990 30080 20070 30100
rect 19990 30040 20010 30080
rect 20050 30040 20070 30080
rect 19990 30020 20070 30040
rect 19930 29960 20010 29990
rect 19870 29900 19950 29930
rect 19750 29010 19830 29040
rect 19750 28870 19780 29010
rect 19810 28960 19890 28980
rect 19810 28920 19830 28960
rect 19870 28920 19890 28960
rect 19810 28900 19890 28920
rect 19750 28840 19830 28870
rect 19690 28780 19770 28810
rect 19740 25170 19770 28780
rect 19610 25140 19770 25170
rect 19610 24960 19640 25140
rect 19670 25060 19770 25080
rect 19670 25020 19690 25060
rect 19730 25020 19770 25060
rect 19670 25000 19770 25020
rect 19550 24940 19640 24960
rect 19550 24930 19580 24940
rect 19560 24900 19580 24930
rect 19620 24900 19640 24940
rect 19560 24880 19640 24900
rect 19740 23850 19770 25000
rect 19690 23830 19770 23850
rect 16700 23530 18200 23830
rect 19690 23790 19710 23830
rect 19750 23790 19770 23830
rect 19690 23770 19770 23790
rect 19800 23680 19830 28840
rect 18260 23650 19830 23680
rect 18260 23530 18290 23650
rect 19860 23620 19890 28900
rect 19920 24960 19950 29900
rect 19980 29170 20010 29960
rect 19980 29150 20060 29170
rect 19980 29110 20000 29150
rect 20040 29110 20060 29150
rect 19980 29090 20060 29110
rect 22860 27260 23010 27330
rect 22780 27250 23010 27260
rect 19920 24930 20140 24960
rect 22930 23760 23010 27250
rect 20340 23740 23010 23760
rect 20340 23700 20360 23740
rect 20400 23700 23010 23740
rect 20340 23680 20420 23700
rect 18320 23590 19890 23620
rect 19990 23620 21820 23650
rect 18320 23530 18350 23590
rect 16640 17830 16700 17890
rect 18420 17770 18480 17830
rect 16640 17710 18480 17770
rect 19990 17630 20050 23620
rect 20090 23570 20170 23590
rect 20090 23530 20110 23570
rect 20150 23530 20170 23570
rect 21790 23530 21820 23620
rect 22930 23530 23010 23700
rect 20090 23510 20170 23530
rect 16640 17570 20050 17630
rect 20110 17510 20170 23510
rect 16640 17450 20170 17510
<< via1 >>
rect 3640 32340 3740 32860
rect 4500 31400 4560 33760
rect 4940 32340 5040 32860
rect 6240 32340 6340 32860
rect 7540 32340 7640 32860
rect 8840 32340 8940 32860
rect 3640 29710 3740 30230
rect 4940 29710 5040 30230
rect 6240 29710 6340 30230
rect 7540 29710 7640 30230
rect 8840 29710 8940 30230
rect 16780 30140 17180 30420
rect 19100 30140 19500 30420
rect 16780 29270 17180 29850
rect 19100 29270 19500 29850
rect 19780 31840 19860 31920
rect 20270 34310 20350 34390
rect 20690 34310 20770 34390
rect 20820 31900 20900 31920
rect 20820 31860 20840 31900
rect 20840 31860 20880 31900
rect 20880 31860 20900 31900
rect 20820 31840 20900 31860
rect 20480 31820 20560 31830
rect 20480 31760 20490 31820
rect 20490 31760 20550 31820
rect 20550 31760 20560 31820
rect 20480 31750 20560 31760
rect 3640 27080 3740 27600
rect 4940 27080 5040 27600
rect 6240 27080 6340 27600
rect 7540 27080 7640 27600
rect 8840 27080 8940 27600
rect 16780 27260 17180 28840
rect 19100 27260 19500 28840
rect 20140 30140 20540 30420
rect 22460 30140 22860 30420
rect 3640 24450 3740 24970
rect 4940 24450 5040 24970
rect 6240 24450 6340 24970
rect 7540 24450 7640 24970
rect 8840 24450 8940 24970
rect 16780 23840 17180 24420
rect 19100 23840 19500 24420
rect 20140 29270 20540 29850
rect 22460 29270 22860 29850
rect 20140 27260 20540 28840
rect 22460 27260 22860 28840
rect 20140 23840 20540 24420
rect 22460 23840 22860 24420
rect 16710 22860 17290 23520
rect 19330 22860 19910 23520
rect 3640 21820 3740 22340
rect 4940 21820 5040 22340
rect 6240 21820 6340 22340
rect 7540 21820 7640 22340
rect 8840 21820 8940 22340
rect 3640 19190 3740 19710
rect 4940 19190 5040 19710
rect 6240 19190 6340 19710
rect 7540 19190 7640 19710
rect 8840 19190 8940 19710
rect 10100 18080 10160 20440
rect 10920 18980 11020 19500
rect 16710 18680 17290 19340
rect 19330 18680 19910 19340
rect 20240 22860 20820 23520
rect 22860 22860 23440 23520
rect 20240 18680 20820 19340
rect 22860 18680 23440 19340
<< metal2 >>
rect 20260 34390 20360 34400
rect 20260 34310 20270 34390
rect 20350 34310 20360 34390
rect 20260 34300 20360 34310
rect 20680 34390 20780 34400
rect 20680 34310 20690 34390
rect 20770 34310 20780 34390
rect 20680 34300 20780 34310
rect 3000 33760 16660 34270
rect 3000 32860 4500 33760
rect 3000 32340 3640 32860
rect 3740 32340 4500 32860
rect 3000 32010 4500 32340
rect 4560 32860 16660 33760
rect 4560 32340 4940 32860
rect 5040 32340 6240 32860
rect 6340 32340 7540 32860
rect 7640 32340 8840 32860
rect 8940 32340 16660 32860
rect 4560 32010 16660 32340
rect 3000 31950 3230 32010
rect 16510 31950 16660 32010
rect 3000 31400 4500 31950
rect 4560 31400 16660 31950
rect 19770 31920 19870 31930
rect 19770 31840 19780 31920
rect 19860 31840 19870 31920
rect 20810 31920 20910 31930
rect 20810 31840 20820 31920
rect 20900 31840 20910 31920
rect 19770 31830 19870 31840
rect 20470 31830 20570 31840
rect 20810 31830 20910 31840
rect 20470 31750 20480 31830
rect 20560 31750 20570 31830
rect 20470 31740 20570 31750
rect 3000 30430 16660 31400
rect 3000 30420 22870 30430
rect 3000 30230 16780 30420
rect 3000 29710 3640 30230
rect 3740 29710 4940 30230
rect 5040 29710 6240 30230
rect 6340 29710 7540 30230
rect 7640 29710 8840 30230
rect 8940 30140 16780 30230
rect 17180 30140 19100 30420
rect 19500 30140 20140 30420
rect 20540 30140 22460 30420
rect 22860 30140 22870 30420
rect 8940 29850 22870 30140
rect 8940 29710 16780 29850
rect 3000 29590 16780 29710
rect 3000 29530 3230 29590
rect 16510 29530 16780 29590
rect 3000 29270 16780 29530
rect 17180 29270 19100 29850
rect 19500 29270 20140 29850
rect 20540 29270 22460 29850
rect 22860 29270 22870 29850
rect 3000 29030 22870 29270
rect 3000 27600 16580 29030
rect 3000 27080 3640 27600
rect 3740 27080 4940 27600
rect 5040 27080 6240 27600
rect 6340 27080 7540 27600
rect 7640 27080 8840 27600
rect 8940 27080 16580 27600
rect 3000 25300 16580 27080
rect 16770 28840 23450 28850
rect 16770 27260 16780 28840
rect 17180 27260 19100 28840
rect 19500 27260 20140 28840
rect 20540 27260 22460 28840
rect 22860 27260 23450 28840
rect 16770 25360 23450 27260
rect 3000 24970 22870 25300
rect 3000 24450 3640 24970
rect 3740 24450 4940 24970
rect 5040 24450 6240 24970
rect 6340 24450 7540 24970
rect 7640 24450 8840 24970
rect 8940 24450 22870 24970
rect 3000 24420 22870 24450
rect 3000 23840 16780 24420
rect 17180 23840 19100 24420
rect 19500 23840 20140 24420
rect 20540 23840 22460 24420
rect 22860 23840 22870 24420
rect 3000 23830 22870 23840
rect 3000 23700 16660 23830
rect 20230 23770 21700 23830
rect 3000 23520 18300 23700
rect 20230 23680 20340 23770
rect 20420 23680 21700 23770
rect 20310 23600 21700 23680
rect 3000 22860 16710 23520
rect 17290 22860 18300 23520
rect 3000 22340 18300 22860
rect 3000 21820 3640 22340
rect 3740 21820 4940 22340
rect 5040 21820 6240 22340
rect 6340 21820 7540 22340
rect 7640 21820 8840 22340
rect 8940 21820 18300 22340
rect 3000 20440 18300 21820
rect 3000 19710 10100 20440
rect 3000 19190 3640 19710
rect 3740 19190 4940 19710
rect 5040 19190 6240 19710
rect 6340 19190 7540 19710
rect 7640 19190 8840 19710
rect 8940 19190 10100 19710
rect 3000 18080 10100 19190
rect 10160 19500 18300 20440
rect 10160 18980 10920 19500
rect 11020 19340 18300 19500
rect 11020 18980 16710 19340
rect 10160 18680 16710 18980
rect 17290 18680 18300 19340
rect 10160 18080 18300 18680
rect 3000 17690 18300 18080
rect 19320 23520 19920 23530
rect 19320 22860 19330 23520
rect 19910 22860 19920 23520
rect 19320 19340 19920 22860
rect 19320 18680 19330 19340
rect 19910 18680 19920 19340
rect 19320 18470 19920 18680
rect 20230 23520 21700 23600
rect 22930 23530 23450 25360
rect 20230 22860 20240 23520
rect 20820 22860 21700 23520
rect 20230 19340 21700 22860
rect 20230 18680 20240 19340
rect 20820 18680 21700 19340
rect 20230 18670 21700 18680
rect 22850 23520 23450 23530
rect 22850 22860 22860 23520
rect 23440 22860 23450 23520
rect 22850 19340 23450 22860
rect 22850 18680 22860 19340
rect 23440 18680 23450 19340
rect 22850 18470 23450 18680
rect 19320 17870 23450 18470
<< via2 >>
rect 20270 34310 20350 34390
rect 20690 34310 20770 34390
rect 3230 31950 4500 32010
rect 4500 31950 4560 32010
rect 4560 31950 16510 32010
rect 19780 31840 19860 31920
rect 20820 31840 20900 31920
rect 20480 31750 20560 31830
rect 3230 29530 16510 29590
<< metal3 >>
rect 18100 34390 22940 34740
rect 18100 34310 20270 34390
rect 20350 34310 20690 34390
rect 20770 34310 22940 34390
rect 18100 34070 22940 34310
rect 3190 32010 23250 34070
rect 3190 31950 3230 32010
rect 16510 31950 16550 32010
rect 3190 31940 16550 31950
rect 19770 31920 19870 31930
rect 19770 31840 19780 31920
rect 19860 31840 19870 31920
rect 20810 31920 20910 31930
rect 20810 31840 20820 31920
rect 20900 31840 20910 31920
rect 19770 31830 19870 31840
rect 20470 31830 20570 31840
rect 20810 31830 20910 31840
rect 20470 31750 20480 31830
rect 20560 31750 20570 31830
rect 3190 29690 23250 31750
rect 3190 29590 16550 29600
rect 3190 29530 3230 29590
rect 16510 29530 16550 29590
rect 3190 17470 23250 29530
<< via3 >>
rect 20270 34310 20350 34390
rect 20690 34310 20770 34390
rect 19780 31840 19860 31920
rect 20820 31840 20900 31920
<< mimcap >>
rect 18130 34610 20130 34710
rect 18130 34310 18630 34610
rect 19630 34310 20130 34610
rect 18130 34210 20130 34310
rect 20910 34610 22910 34710
rect 20910 34310 21410 34610
rect 22410 34310 22910 34610
rect 20910 34210 22910 34310
rect 3220 33540 23220 34040
rect 3220 32540 18220 33540
rect 20220 32540 23220 33540
rect 3220 32040 23220 32540
rect 3220 31210 23220 31720
rect 3220 30210 18220 31210
rect 20220 30210 23220 31210
rect 3220 29720 23220 30210
rect 3220 26540 23220 29500
rect 3220 24540 18220 26540
rect 20220 24540 23220 26540
rect 3220 17500 23220 24540
<< mimcapcontact >>
rect 18630 34310 19630 34610
rect 21410 34310 22410 34610
rect 18220 32540 20220 33540
rect 18220 30210 20220 31210
rect 18220 24540 20220 26540
<< metal4 >>
rect 18620 34610 19640 34620
rect 18620 34310 18630 34610
rect 19630 34400 19640 34610
rect 21400 34610 22420 34620
rect 21400 34400 21410 34610
rect 19630 34390 20360 34400
rect 19630 34310 20270 34390
rect 20350 34310 20360 34390
rect 18620 34300 20360 34310
rect 20680 34390 21410 34400
rect 20680 34310 20690 34390
rect 20770 34310 21410 34390
rect 22410 34310 22420 34610
rect 20680 34300 22420 34310
rect 18210 33540 20230 33550
rect 18210 32540 18220 33540
rect 20220 32540 20230 33540
rect 18210 32530 20230 32540
rect 19770 31920 19870 32530
rect 19770 31840 19780 31920
rect 19860 31840 19870 31920
rect 19770 31830 19870 31840
rect 20810 31920 20910 31930
rect 20810 31840 20820 31920
rect 20900 31840 20910 31920
rect 20810 31220 20910 31840
rect 18210 31210 20910 31220
rect 18210 30210 18220 31210
rect 20220 31120 20910 31210
rect 20220 30210 20230 31120
rect 18210 30200 20230 30210
rect 20130 26550 20230 30200
rect 20810 26550 20910 30650
rect 18210 26540 20910 26550
rect 18210 24540 18220 26540
rect 20220 26450 20910 26540
rect 20220 24540 20230 26450
rect 18210 24530 20230 24540
use 4_bit_binary_decoder  4_bit_binary_decoder_0
timestamp 1702679905
transform 1 0 2780 0 1 34820
box -73 -54 3780 971
use bias  bias_0
timestamp 1697165931
transform 0 1 16780 1 0 19350
box -1560 -150 4220 3210
use bias  bias_1
timestamp 1697165931
transform 0 1 20310 1 0 19350
box -1560 -150 4220 3210
use current_steering_dac  current_steering_dac_0
timestamp 1702726065
transform 1 0 10080 0 1 18030
box -7300 -580 6560 16450
use opamp_balanced  opamp_balanced_0
timestamp 1702677968
transform -1 0 19410 0 1 24570
box -140 -870 2770 6050
use opamp_balanced  opamp_balanced_1
timestamp 1702677968
transform 1 0 20230 0 1 24570
box -140 -870 2770 6050
use switched_capacitor_transmission_gate  switched_capacitor_transmission_gate_0
timestamp 1702761464
transform 1 0 20130 0 1 30770
box -40 -30 400 3420
use switched_capacitor_transmission_gate  switched_capacitor_transmission_gate_1
timestamp 1702761464
transform 1 0 20550 0 1 30770
box -40 -30 400 3420
<< labels >>
flabel metal1 19990 35750 19990 35750 1 FreeSans 800 0 0 0 Vref
flabel locali 23520 30720 23520 30720 3 FreeSans 800 0 0 0 Vout
flabel locali 21900 17450 21900 17450 5 FreeSans 800 0 0 0 Ibdac
flabel locali 18370 17450 18370 17450 5 FreeSans 800 0 0 0 Ibfilter
<< end >>
