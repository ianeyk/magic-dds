magic
tech sky130A
magscale 1 2
timestamp 1702722287
<< error_p >>
rect 3728 19710 3740 19712
rect 5028 19710 5040 19712
rect 6328 19710 6340 19712
rect 7628 19710 7640 19712
rect 8928 19710 8940 19712
rect 3750 19688 3752 19700
rect 5050 19688 5052 19700
rect 6350 19688 6352 19700
rect 7650 19688 7652 19700
rect 8950 19688 8952 19700
rect 10908 18990 10910 19002
rect 12208 18990 12210 19002
rect 13508 18990 13510 19002
rect 14808 18990 14810 19002
rect 10920 18978 10932 18980
rect 12220 18978 12232 18980
rect 13520 18978 13532 18980
rect 14820 18978 14832 18980
<< error_s >>
rect 3728 32860 3740 32862
rect 5028 32860 5040 32862
rect 6328 32860 6340 32862
rect 7628 32860 7640 32862
rect 8928 32860 8940 32862
rect 3750 32838 3752 32850
rect 5050 32838 5052 32850
rect 6350 32838 6352 32850
rect 7650 32838 7652 32850
rect 8950 32838 8952 32850
rect 10908 32140 10910 32152
rect 12208 32140 12210 32152
rect 13508 32140 13510 32152
rect 14808 32140 14810 32152
rect 16108 32140 16110 32152
rect 10920 32128 10932 32130
rect 12220 32128 12232 32130
rect 13520 32128 13532 32130
rect 14820 32128 14832 32130
rect 16120 32128 16132 32130
rect 3728 30230 3740 30232
rect 3750 30208 3752 30220
rect 16108 29510 16110 29522
rect 16120 29498 16132 29500
rect 9810 28630 9814 28650
rect 9776 28610 9780 28630
rect 3728 27600 3740 27602
rect 3750 27578 3752 27590
rect 16108 26880 16110 26892
rect 16120 26868 16132 26870
rect 3728 24970 3740 24972
rect 3750 24948 3752 24960
rect 16108 24250 16110 24262
rect 16120 24238 16132 24240
rect 3728 22340 3740 22342
rect 3750 22318 3752 22330
rect 16108 21620 16110 21632
rect 16120 21608 16132 21610
rect 16108 18990 16110 19002
rect 16120 18978 16132 18980
<< locali >>
rect 2780 34680 2820 34820
rect 3460 34680 3500 34820
rect 2780 34660 2960 34680
rect 2780 34640 2900 34660
rect 2880 34620 2900 34640
rect 2940 34620 2960 34660
rect 2880 34600 2960 34620
rect 2920 34480 2960 34600
rect 3000 34640 3500 34680
rect 3000 34480 3040 34640
rect 3880 34600 3920 34820
rect 3080 34560 3920 34600
rect 3080 34480 3120 34560
rect 4140 34520 4180 34820
rect 4670 34740 4710 34820
rect 5350 34740 5390 34820
rect 5770 34740 5810 34820
rect 5900 34780 6070 34820
rect 4670 34720 4750 34740
rect 4670 34680 4690 34720
rect 4730 34680 4750 34720
rect 4670 34660 4750 34680
rect 5350 34720 5430 34740
rect 5350 34680 5370 34720
rect 5410 34680 5430 34720
rect 5350 34660 5430 34680
rect 5770 34720 5850 34740
rect 5770 34680 5790 34720
rect 5830 34680 5850 34720
rect 5770 34660 5850 34680
rect 3160 34480 4180 34520
rect 5900 34480 5940 34780
rect 5980 34720 6060 34740
rect 5980 34680 6000 34720
rect 6040 34680 6060 34720
rect 5980 34660 6060 34680
rect 5980 34480 6020 34660
rect 6100 34640 6180 34660
rect 6100 34620 6120 34640
rect 6060 34600 6120 34620
rect 6160 34600 6180 34640
rect 6060 34580 6180 34600
rect 6220 34580 6300 34600
rect 6060 34480 6100 34580
rect 6220 34540 6240 34580
rect 6280 34540 6300 34580
rect 6220 34520 6300 34540
rect 6140 34480 6260 34520
rect 19510 33900 19940 33920
rect 19510 33880 19880 33900
rect 19860 33860 19880 33880
rect 19920 33860 19940 33900
rect 19860 33840 19940 33860
rect 19500 33260 20290 33280
rect 19500 33220 20230 33260
rect 20270 33220 20290 33260
rect 19500 33200 20290 33220
rect 19510 33090 19770 33110
rect 19510 33070 19710 33090
rect 19690 33050 19710 33070
rect 19750 33050 19770 33090
rect 19690 33030 19770 33050
rect 19570 31880 19650 31900
rect 19570 31840 19590 31880
rect 19630 31860 19650 31880
rect 19630 31840 19960 31860
rect 19570 31820 19960 31840
rect 19510 31420 19710 31440
rect 19510 31400 19650 31420
rect 19630 31380 19650 31400
rect 19690 31380 19710 31420
rect 19630 31360 19710 31380
rect 19510 30600 19880 30620
rect 19510 30580 19820 30600
rect 19800 30560 19820 30580
rect 19860 30560 19880 30600
rect 19800 30540 19880 30560
rect 19920 30060 19960 31820
rect 19510 30020 19960 30060
rect 20000 30580 20350 30620
rect 20000 29980 20040 30580
rect 19800 29960 20040 29980
rect 19800 29920 19820 29960
rect 19860 29940 20040 29960
rect 19860 29920 19880 29940
rect 19800 29900 19880 29920
rect 19500 29770 20360 29850
rect 19510 29090 19970 29130
rect 20170 29090 20350 29130
rect 19510 28960 20350 28980
rect 19510 28940 19880 28960
rect 19860 28920 19880 28940
rect 19920 28940 20350 28960
rect 19920 28920 19940 28940
rect 19860 28900 19940 28920
rect 19500 27320 20360 27340
rect 19500 27280 20230 27320
rect 20270 27280 20360 27320
rect 19500 27260 20360 27280
rect 19510 27150 20350 27170
rect 19510 27130 19710 27150
rect 19670 27110 19710 27130
rect 19750 27130 20350 27150
rect 19750 27110 19770 27130
rect 19670 27090 19770 27110
rect 19550 25180 19630 25200
rect 19550 25140 19570 25180
rect 19610 25140 19630 25180
rect 19550 25120 19630 25140
rect 19550 24500 19590 25120
rect 19670 25080 19710 27090
rect 19670 25060 19750 25080
rect 19670 25020 19690 25060
rect 19730 25020 19750 25060
rect 19670 25000 19750 25020
rect 19630 24940 19930 24960
rect 19630 24900 19650 24940
rect 19690 24920 19930 24940
rect 19690 24900 19710 24920
rect 19630 24880 19710 24900
rect 19510 24460 20350 24500
rect 19550 23930 19590 24460
rect 19550 23910 20170 23930
rect 19550 23890 20110 23910
rect 19550 23680 19590 23890
rect 20090 23870 20110 23890
rect 20150 23870 20170 23910
rect 20090 23850 20170 23870
rect 18200 23640 19590 23680
rect 19670 23830 19770 23850
rect 19670 23790 19710 23830
rect 19750 23790 19770 23830
rect 19670 23770 19770 23790
rect 18200 23530 18240 23640
rect 19670 23600 19710 23770
rect 19750 23710 19830 23730
rect 19750 23670 19770 23710
rect 19810 23690 19830 23710
rect 19810 23670 20050 23690
rect 19750 23650 19990 23670
rect 19970 23630 19990 23650
rect 20030 23630 20050 23670
rect 19970 23610 20050 23630
rect 18380 23560 19710 23600
rect 18380 23530 18420 23560
rect 19890 23500 20310 23520
rect 19890 23460 20250 23500
rect 20290 23460 20310 23500
rect 19890 23440 20310 23460
<< viali >>
rect 2900 34620 2940 34660
rect 4690 34680 4730 34720
rect 5370 34680 5410 34720
rect 5790 34680 5830 34720
rect 6000 34680 6040 34720
rect 6120 34600 6160 34640
rect 6240 34540 6280 34580
rect 19880 33860 19920 33900
rect 20230 33220 20270 33260
rect 19710 33050 19750 33090
rect 19590 31840 19630 31880
rect 19650 31380 19690 31420
rect 19820 30560 19860 30600
rect 19820 29920 19860 29960
rect 19880 28920 19920 28960
rect 20230 27280 20270 27320
rect 19710 27110 19750 27150
rect 19570 25140 19610 25180
rect 19690 25020 19730 25060
rect 19650 24900 19690 24940
rect 20110 23870 20150 23910
rect 19710 23790 19750 23830
rect 19770 23670 19810 23710
rect 19990 23630 20030 23670
rect 20250 23460 20290 23500
<< metal1 >>
rect 2880 34660 2960 34680
rect 2880 34620 2900 34660
rect 2940 34620 3080 34660
rect 2880 34600 3080 34620
rect 3020 34480 3080 34600
rect 3160 34480 3220 34850
rect 4670 34720 4750 34740
rect 4670 34680 4690 34720
rect 4730 34680 4750 34720
rect 4670 34660 4750 34680
rect 5350 34720 5430 34740
rect 5350 34680 5370 34720
rect 5410 34680 5430 34720
rect 5350 34660 5430 34680
rect 5770 34720 5850 34740
rect 5770 34680 5790 34720
rect 5830 34690 5850 34720
rect 5980 34720 6060 34740
rect 5980 34690 6000 34720
rect 5830 34680 6000 34690
rect 6040 34680 6060 34720
rect 5770 34660 6060 34680
rect 4720 34550 4750 34660
rect 5400 34610 5430 34660
rect 6100 34640 6180 34660
rect 6100 34610 6120 34640
rect 5400 34600 6120 34610
rect 6160 34600 6180 34640
rect 5400 34580 6180 34600
rect 6220 34580 6300 34600
rect 6220 34550 6240 34580
rect 4720 34540 6240 34550
rect 6280 34540 6300 34580
rect 4720 34520 6300 34540
rect 16640 34400 17770 34460
rect 16640 34280 17380 34340
rect 17320 33980 17380 34280
rect 17710 33900 17770 34400
rect 19860 33900 19940 33920
rect 19860 33860 19880 33900
rect 19920 33860 19940 33900
rect 19860 33840 19940 33860
rect 19690 33090 19770 33110
rect 19690 33050 19710 33090
rect 19750 33050 19770 33090
rect 19690 33030 19770 33050
rect 19550 31880 19650 31900
rect 19550 31870 19590 31880
rect 19570 31840 19590 31870
rect 19630 31840 19650 31880
rect 19570 31820 19650 31840
rect 19630 31420 19710 31440
rect 19630 31380 19650 31420
rect 19690 31380 19710 31420
rect 19630 31360 19710 31380
rect 16640 30770 16770 30830
rect 19630 25200 19660 31360
rect 19740 27170 19770 33030
rect 19690 27150 19770 27170
rect 19690 27110 19710 27150
rect 19750 27110 19770 27150
rect 19690 27090 19770 27110
rect 19800 30600 19880 30620
rect 19800 30560 19820 30600
rect 19860 30560 19880 30600
rect 19800 30540 19880 30560
rect 19800 29980 19830 30540
rect 19800 29960 19880 29980
rect 19800 29920 19820 29960
rect 19860 29920 19880 29960
rect 19800 29900 19880 29920
rect 19550 25180 19660 25200
rect 19550 25140 19570 25180
rect 19610 25140 19660 25180
rect 19550 25120 19660 25140
rect 19670 25060 19770 25080
rect 19670 25020 19690 25060
rect 19730 25020 19770 25060
rect 19670 25000 19770 25020
rect 19550 24940 19710 24960
rect 19550 24930 19650 24940
rect 19630 24900 19650 24930
rect 19690 24900 19710 24940
rect 19630 24880 19710 24900
rect 19740 23850 19770 25000
rect 19690 23830 19770 23850
rect 16700 23530 18200 23830
rect 19690 23790 19710 23830
rect 19750 23790 19770 23830
rect 19690 23770 19770 23790
rect 19800 23730 19830 29900
rect 19910 28980 19940 33840
rect 20210 33260 20290 33280
rect 20210 33220 20230 33260
rect 20270 33220 20290 33260
rect 20210 33200 20290 33220
rect 19750 23710 19830 23730
rect 19750 23680 19770 23710
rect 18260 23670 19770 23680
rect 19810 23670 19830 23710
rect 18260 23650 19830 23670
rect 19860 28960 19940 28980
rect 19860 28920 19880 28960
rect 19920 28920 19940 28960
rect 19860 28900 19940 28920
rect 18260 23530 18290 23650
rect 19860 23620 19890 28900
rect 20230 27340 20290 33200
rect 20210 27320 20290 27340
rect 20210 27280 20230 27320
rect 20270 27280 20290 27320
rect 20210 27260 20290 27280
rect 20230 25080 20290 27260
rect 20220 24990 20290 25080
rect 20220 24900 20280 24990
rect 20220 24810 20290 24900
rect 20090 23910 20170 23930
rect 20090 23870 20110 23910
rect 20150 23870 20170 23910
rect 20090 23850 20170 23870
rect 18320 23590 19890 23620
rect 19970 23670 20050 23690
rect 19970 23630 19990 23670
rect 20030 23630 20050 23670
rect 19970 23610 20050 23630
rect 18320 23530 18350 23590
rect 16640 17830 16700 17890
rect 18420 17770 18480 17830
rect 16640 17710 18480 17770
rect 19990 17630 20050 23610
rect 16640 17570 20050 17630
rect 20110 17510 20170 23850
rect 20230 23520 20290 24810
rect 20230 23500 20310 23520
rect 20230 23460 20250 23500
rect 20290 23460 20310 23500
rect 20230 23440 20310 23460
rect 16640 17450 20170 17510
use 4_bit_binary_decoder  4_bit_binary_decoder_0
timestamp 1702679905
transform 1 0 2780 0 1 34820
box -73 -54 3780 971
use bias  bias_0
timestamp 1697165931
transform 0 1 16780 1 0 19350
box -1560 -150 4220 3210
use current_difference_balanced  current_difference_balanced_0
timestamp 1702677849
transform -1 0 19410 0 1 31510
box -140 -870 2680 2500
use current_steering_dac  current_steering_dac_0
timestamp 1702722181
transform 1 0 10080 0 1 18030
box -7300 -580 6560 16450
use opamp_balanced  opamp_balanced_0
timestamp 1702677968
transform -1 0 19410 0 1 24570
box -140 -870 2770 6050
use opamp_balanced  opamp_balanced_1
timestamp 1702677968
transform 1 0 20450 0 1 24570
box -140 -870 2770 6050
use switched_capacitor_transmission_gate  switched_capacitor_transmission_gate_0
timestamp 1702721627
transform 1 0 20690 0 1 30930
box -40 -110 400 3420
<< end >>
