magic
tech sky130A
magscale 1 2
timestamp 1702759971
<< error_s >>
rect 20770 31640 20944 34120
<< xpolycontact >>
rect 16780 33480 16920 33920
rect 16780 30740 16920 31180
rect 17170 33480 17310 33920
rect 17170 30740 17310 31180
rect 17560 33480 17700 33920
rect 17560 30740 17700 31180
rect 17950 33480 18090 33920
rect 17950 30740 18090 31180
rect 18340 33480 18480 33920
rect 18340 30740 18480 31180
rect 18730 33480 18870 33920
rect 18730 30740 18870 31180
<< xpolyres >>
rect 16780 31180 16920 33480
rect 17170 31180 17310 33480
rect 17560 31180 17700 33480
rect 17950 31180 18090 33480
rect 18340 31180 18480 33480
rect 18730 31180 18870 33480
<< locali >>
rect 2780 34680 2820 34820
rect 3460 34680 3500 34820
rect 2780 34660 2960 34680
rect 2780 34640 2900 34660
rect 2880 34620 2900 34640
rect 2940 34620 2960 34660
rect 2880 34600 2960 34620
rect 2920 34480 2960 34600
rect 3000 34640 3500 34680
rect 3000 34480 3040 34640
rect 3880 34600 3920 34820
rect 3080 34560 3920 34600
rect 3080 34480 3120 34560
rect 4140 34520 4180 34820
rect 4670 34740 4710 34820
rect 5350 34740 5390 34820
rect 5770 34740 5810 34820
rect 5900 34780 6070 34820
rect 4670 34720 4750 34740
rect 4670 34680 4690 34720
rect 4730 34680 4750 34720
rect 4670 34660 4750 34680
rect 5350 34720 5430 34740
rect 5350 34680 5370 34720
rect 5410 34680 5430 34720
rect 5350 34660 5430 34680
rect 5770 34720 5850 34740
rect 5770 34680 5790 34720
rect 5830 34680 5850 34720
rect 5770 34660 5850 34680
rect 3160 34480 4180 34520
rect 5900 34480 5940 34780
rect 5980 34720 6060 34740
rect 5980 34680 6000 34720
rect 6040 34680 6060 34720
rect 5980 34660 6060 34680
rect 5980 34480 6020 34660
rect 6100 34640 6180 34660
rect 6100 34620 6120 34640
rect 6060 34600 6120 34620
rect 6160 34600 6180 34640
rect 6060 34580 6180 34600
rect 6220 34580 6300 34600
rect 6060 34480 6100 34580
rect 6220 34540 6240 34580
rect 6280 34540 6300 34580
rect 6220 34520 6300 34540
rect 6140 34480 6260 34520
rect 17170 34460 17250 34480
rect 17170 34420 17190 34460
rect 17230 34420 17250 34460
rect 16780 34320 16860 34340
rect 16780 34280 16800 34320
rect 16840 34280 16860 34320
rect 16780 33920 16860 34280
rect 17170 33920 17250 34420
rect 18010 34000 18810 34080
rect 18010 33920 18090 34000
rect 18730 33920 18810 34000
rect 17620 33400 17700 33480
rect 18340 33400 18420 33480
rect 17620 33320 18420 33400
rect 16840 31270 17640 31340
rect 16840 31180 16920 31270
rect 17560 31180 17640 31270
rect 18400 31320 19820 31340
rect 18400 31280 19760 31320
rect 19800 31280 19820 31320
rect 18400 31260 19820 31280
rect 18400 31180 18480 31260
rect 17230 30650 17310 30740
rect 17950 30650 18030 30740
rect 17230 30580 18030 30650
rect 19510 30600 20350 30620
rect 19510 30580 19820 30600
rect 19800 30560 19820 30580
rect 19860 30580 20350 30600
rect 19860 30560 19880 30580
rect 19800 30540 19880 30560
rect 19570 30080 19650 30100
rect 19570 30060 19590 30080
rect 19510 30040 19590 30060
rect 19630 30040 19650 30080
rect 19510 30020 19650 30040
rect 19990 30080 20070 30100
rect 19990 30040 20010 30080
rect 20050 30060 20070 30080
rect 20050 30040 20130 30060
rect 19990 30020 20130 30040
rect 19500 29770 20360 29850
rect 19630 29190 19710 29210
rect 19630 29150 19650 29190
rect 19690 29150 19710 29190
rect 19630 29130 19710 29150
rect 19980 29150 20060 29170
rect 19510 29090 19670 29130
rect 19980 29110 20000 29150
rect 20040 29130 20060 29150
rect 20040 29110 20130 29130
rect 19980 29090 20130 29110
rect 20170 29090 20350 29130
rect 19510 28960 20350 28980
rect 19510 28940 19830 28960
rect 19810 28920 19830 28940
rect 19870 28940 20350 28960
rect 19870 28920 19890 28940
rect 19810 28900 19890 28920
rect 19500 27260 20360 27340
rect 19510 27130 20350 27170
rect 19670 25080 19710 27130
rect 19670 25060 19750 25080
rect 19670 25020 19690 25060
rect 19730 25020 19750 25060
rect 19670 25000 19750 25020
rect 19560 24940 19640 24960
rect 19560 24900 19580 24940
rect 19620 24900 19640 24940
rect 19560 24880 19640 24900
rect 19510 24460 20350 24500
rect 19550 23930 19590 24460
rect 19550 23890 19960 23930
rect 19550 23680 19590 23890
rect 18200 23640 19590 23680
rect 19670 23830 19770 23850
rect 19670 23790 19710 23830
rect 19750 23790 19770 23830
rect 19670 23770 19770 23790
rect 19920 23770 19960 23890
rect 18200 23530 18240 23640
rect 19670 23600 19710 23770
rect 19920 23750 20000 23770
rect 19750 23710 19830 23730
rect 19750 23670 19770 23710
rect 19810 23670 19830 23710
rect 19920 23710 19940 23750
rect 19980 23710 20000 23750
rect 19920 23690 20000 23710
rect 19750 23650 19830 23670
rect 19790 23630 20050 23650
rect 19790 23610 19990 23630
rect 18380 23560 19710 23600
rect 19970 23590 19990 23610
rect 20030 23590 20050 23630
rect 19970 23570 20050 23590
rect 18380 23530 18420 23560
rect 19890 23500 20310 23520
rect 19890 23460 20250 23500
rect 20290 23460 20310 23500
rect 19890 23440 20310 23460
<< viali >>
rect 2900 34620 2940 34660
rect 4690 34680 4730 34720
rect 5370 34680 5410 34720
rect 5790 34680 5830 34720
rect 6000 34680 6040 34720
rect 6120 34600 6160 34640
rect 6240 34540 6280 34580
rect 17190 34420 17230 34460
rect 16800 34280 16840 34320
rect 19760 31280 19800 31320
rect 19820 30560 19860 30600
rect 19590 30040 19630 30080
rect 20010 30040 20050 30080
rect 19650 29150 19690 29190
rect 20000 29110 20040 29150
rect 19830 28920 19870 28960
rect 19690 25020 19730 25060
rect 19580 24900 19620 24940
rect 19710 23790 19750 23830
rect 19770 23670 19810 23710
rect 19940 23710 19980 23750
rect 19990 23590 20030 23630
rect 20250 23460 20290 23500
<< metal1 >>
rect 2880 34660 2960 34680
rect 2880 34620 2900 34660
rect 2940 34620 3080 34660
rect 2880 34600 3080 34620
rect 3020 34480 3080 34600
rect 3160 34480 3220 34850
rect 4670 34720 4750 34740
rect 4670 34680 4690 34720
rect 4730 34680 4750 34720
rect 4670 34660 4750 34680
rect 5350 34720 5430 34740
rect 5350 34680 5370 34720
rect 5410 34680 5430 34720
rect 5350 34660 5430 34680
rect 5770 34720 5850 34740
rect 5770 34680 5790 34720
rect 5830 34690 5850 34720
rect 5980 34720 6060 34740
rect 5980 34690 6000 34720
rect 5830 34680 6000 34690
rect 6040 34680 6060 34720
rect 5770 34660 6060 34680
rect 4720 34550 4750 34660
rect 5400 34610 5430 34660
rect 6100 34640 6180 34660
rect 6100 34610 6120 34640
rect 5400 34600 6120 34610
rect 6160 34600 6180 34640
rect 5400 34580 6180 34600
rect 6220 34580 6300 34600
rect 6220 34550 6240 34580
rect 4720 34540 6240 34550
rect 6280 34540 6300 34580
rect 4720 34520 6300 34540
rect 17170 34460 17250 34480
rect 16640 34420 17190 34460
rect 17230 34420 19710 34460
rect 16640 34400 19710 34420
rect 16640 34320 19600 34340
rect 16640 34280 16800 34320
rect 16840 34280 19600 34320
rect 16780 34260 16860 34280
rect 19570 30100 19600 34280
rect 19570 30080 19650 30100
rect 19570 30040 19590 30080
rect 19630 30040 19650 30080
rect 19570 30020 19650 30040
rect 19680 29210 19710 34400
rect 19630 29190 19710 29210
rect 19630 29150 19650 29190
rect 19690 29150 19710 29190
rect 19630 29130 19710 29150
rect 19740 31340 19770 34810
rect 19740 31320 19820 31340
rect 19740 31280 19760 31320
rect 19800 31280 19820 31320
rect 19740 31260 19820 31280
rect 19740 29100 19770 31260
rect 19690 29070 19770 29100
rect 19800 30600 19880 30620
rect 19800 30560 19820 30600
rect 19860 30560 19880 30600
rect 19800 30540 19880 30560
rect 19690 28810 19720 29070
rect 19800 29040 19830 30540
rect 19920 30220 19950 35000
rect 19870 30190 19950 30220
rect 19870 29930 19900 30190
rect 19980 30160 20010 35000
rect 19930 30130 20010 30160
rect 19930 29990 19960 30130
rect 20040 30100 20070 35000
rect 19990 30080 20070 30100
rect 19990 30040 20010 30080
rect 20050 30040 20070 30080
rect 19990 30020 20070 30040
rect 19930 29960 20010 29990
rect 19870 29900 19950 29930
rect 19750 29010 19830 29040
rect 19750 28870 19780 29010
rect 19810 28960 19890 28980
rect 19810 28920 19830 28960
rect 19870 28920 19890 28960
rect 19810 28900 19890 28920
rect 19750 28840 19830 28870
rect 19690 28780 19770 28810
rect 19740 25170 19770 28780
rect 19610 25140 19770 25170
rect 19610 24960 19640 25140
rect 19670 25060 19770 25080
rect 19670 25020 19690 25060
rect 19730 25020 19770 25060
rect 19670 25000 19770 25020
rect 19550 24940 19640 24960
rect 19550 24930 19580 24940
rect 19560 24900 19580 24930
rect 19620 24900 19640 24940
rect 19560 24880 19640 24900
rect 19740 23850 19770 25000
rect 19690 23830 19770 23850
rect 16700 23530 18200 23830
rect 19690 23790 19710 23830
rect 19750 23790 19770 23830
rect 19690 23770 19770 23790
rect 19800 23730 19830 28840
rect 19750 23710 19830 23730
rect 19750 23680 19770 23710
rect 18260 23670 19770 23680
rect 19810 23670 19830 23710
rect 18260 23650 19830 23670
rect 18260 23530 18290 23650
rect 19860 23620 19890 28900
rect 19920 24960 19950 29900
rect 19980 29170 20010 29960
rect 19980 29150 20060 29170
rect 19980 29110 20000 29150
rect 20040 29110 20060 29150
rect 19980 29090 20060 29110
rect 19920 24930 20140 24960
rect 19920 23750 20000 23770
rect 19920 23710 19940 23750
rect 19980 23710 20170 23750
rect 19920 23690 20170 23710
rect 18320 23590 19890 23620
rect 19970 23630 20050 23650
rect 19970 23590 19990 23630
rect 20030 23590 20050 23630
rect 18320 23530 18350 23590
rect 19970 23570 20050 23590
rect 16640 17830 16700 17890
rect 18420 17770 18480 17830
rect 16640 17710 18480 17770
rect 19990 17630 20050 23570
rect 16640 17570 20050 17630
rect 20110 17510 20170 23690
rect 20230 23500 20310 23520
rect 20230 23460 20250 23500
rect 20290 23460 20310 23500
rect 20230 23440 20310 23460
rect 16640 17450 20170 17510
use 4_bit_binary_decoder  4_bit_binary_decoder_0
timestamp 1702679905
transform 1 0 2780 0 1 34820
box -73 -54 3780 971
use bias  bias_0
timestamp 1697165931
transform 0 1 16780 1 0 19350
box -1560 -150 4220 3210
use current_steering_dac  current_steering_dac_0
timestamp 1702726065
transform 1 0 10080 0 1 18030
box -7300 -580 6560 16450
use opamp_balanced  opamp_balanced_0
timestamp 1702677968
transform -1 0 19410 0 1 24570
box -140 -870 2770 6050
use opamp_balanced  opamp_balanced_1
timestamp 1702677968
transform 1 0 20230 0 1 24570
box -140 -870 2770 6050
use switched_capacitor_transmission_gate  switched_capacitor_transmission_gate_0
timestamp 1702744874
transform 1 0 20290 0 1 30770
box -40 -110 400 3420
use switched_capacitor_transmission_gate  switched_capacitor_transmission_gate_1
timestamp 1702744874
transform 1 0 20810 0 1 30770
box -40 -110 400 3420
<< end >>
