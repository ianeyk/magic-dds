magic
tech sky130A
timestamp 1702743177
<< nwell >>
rect -95 180 270 320
<< nmos >>
rect 50 0 65 100
rect 90 0 105 100
rect 130 0 145 100
<< pmos >>
rect 25 200 40 300
rect 90 200 105 300
rect 155 200 170 300
<< ndiff >>
rect 0 85 50 100
rect 0 15 15 85
rect 35 15 50 85
rect 0 0 50 15
rect 65 0 90 100
rect 105 0 130 100
rect 145 85 195 100
rect 145 15 160 85
rect 180 15 195 85
rect 145 0 195 15
<< pdiff >>
rect -25 285 25 300
rect -25 215 -10 285
rect 10 215 25 285
rect -25 200 25 215
rect 40 285 90 300
rect 40 215 55 285
rect 75 215 90 285
rect 40 200 90 215
rect 105 285 155 300
rect 105 215 120 285
rect 140 215 155 285
rect 105 200 155 215
rect 170 280 220 300
rect 170 215 185 280
rect 205 215 220 280
rect 170 200 220 215
<< ndiffc >>
rect 15 15 35 85
rect 160 15 180 85
<< pdiffc >>
rect -10 215 10 285
rect 55 215 75 285
rect 120 215 140 285
rect 185 215 205 280
<< psubdiff >>
rect -50 85 0 100
rect -50 15 -35 85
rect -15 15 0 85
rect -50 0 0 15
<< nsubdiff >>
rect -75 285 -25 300
rect -75 215 -60 285
rect -40 215 -25 285
rect -75 200 -25 215
<< psubdiffcont >>
rect -35 15 -15 85
<< nsubdiffcont >>
rect -60 215 -40 285
<< poly >>
rect 25 300 40 315
rect 90 300 105 315
rect 155 300 170 315
rect 25 165 40 200
rect 25 150 65 165
rect 50 100 65 150
rect 90 100 105 200
rect 155 165 170 200
rect 130 150 170 165
rect 130 100 145 150
rect 50 -15 65 0
rect 90 -15 105 0
rect 130 -15 145 0
<< locali >>
rect -70 285 20 295
rect -70 215 -60 285
rect -40 215 -10 285
rect 10 215 20 285
rect -70 205 20 215
rect 45 285 85 295
rect 45 215 55 285
rect 75 215 85 285
rect 45 205 85 215
rect 110 285 150 295
rect 110 215 120 285
rect 140 215 150 285
rect 110 205 150 215
rect 175 280 215 295
rect 175 215 185 280
rect 205 215 215 280
rect 175 205 215 215
rect 65 155 85 205
rect 175 155 195 205
rect 65 135 195 155
rect 150 95 170 135
rect -45 85 45 95
rect -45 15 -35 85
rect -15 15 15 85
rect 35 15 45 85
rect -45 5 45 15
rect 150 85 190 95
rect 150 15 160 85
rect 180 15 190 85
rect 150 5 190 15
<< viali >>
rect -60 215 -40 285
rect -10 215 10 285
rect 120 215 140 285
<< metal1 >>
rect -70 285 150 295
rect -70 215 -60 285
rect -40 215 -10 285
rect 10 215 120 285
rect 140 215 150 285
rect -70 205 150 215
rect 175 205 215 295
<< labels >>
flabel poly 55 -15 55 -15 1 FreeSans 160 0 0 0 A
port 1 n
flabel poly 95 -15 95 -15 1 FreeSans 160 0 0 0 B
port 2 n
flabel locali 65 295 65 295 5 FreeSans 160 0 0 0 Y
port 3 s
flabel locali -45 50 -45 50 3 FreeSans 160 0 0 0 VN
port 5 e
flabel locali -70 250 -70 250 3 FreeSans 160 0 0 0 VP
port 4 e
flabel poly 135 -15 135 -15 1 FreeSans 160 0 0 0 C
port 6 n
<< end >>
