magic
tech sky130A
magscale 1 2
timestamp 1702591987
<< error_s >>
rect -6352 14830 -6340 14832
rect -5052 14830 -5040 14832
rect -3752 14830 -3740 14832
rect -2452 14830 -2440 14832
rect -1152 14830 -1140 14832
rect -6330 14808 -6328 14820
rect -5030 14808 -5028 14820
rect -3730 14808 -3728 14820
rect -2430 14808 -2428 14820
rect -1130 14808 -1128 14820
rect 828 14110 830 14122
rect 2128 14110 2130 14122
rect 3428 14110 3430 14122
rect 4728 14110 4730 14122
rect 6028 14110 6030 14122
rect 840 14098 852 14100
rect 2140 14098 2152 14100
rect 3440 14098 3452 14100
rect 4740 14098 4752 14100
rect 6040 14098 6052 14100
rect -1152 12200 -1140 12202
rect -1130 12178 -1128 12190
rect 828 11480 830 11492
rect 840 11468 852 11470
rect -270 10600 -266 10620
rect -304 10580 -300 10600
rect -1152 9570 -1140 9572
rect -1130 9548 -1128 9560
rect 828 8850 830 8862
rect 840 8838 852 8840
rect -1152 6940 -1140 6942
rect -1130 6918 -1128 6930
rect 828 6220 830 6232
rect 840 6208 852 6210
rect -1152 4310 -1140 4312
rect -1130 4288 -1128 4300
rect 828 3590 830 3602
rect 840 3578 852 3580
rect -6352 1680 -6340 1682
rect -5052 1680 -5040 1682
rect -3752 1680 -3740 1682
rect -2452 1680 -2440 1682
rect -1152 1680 -1140 1682
rect -6330 1658 -6328 1670
rect -5030 1658 -5028 1670
rect -3730 1658 -3728 1670
rect -2430 1658 -2428 1670
rect -1130 1658 -1128 1670
rect 828 960 830 972
rect 2128 960 2130 972
rect 3428 960 3430 972
rect 4728 960 4730 972
rect 6028 960 6030 972
rect 840 948 852 950
rect 2140 948 2152 950
rect 3440 948 3452 950
rect 4740 948 4752 950
rect 6040 948 6052 950
<< poly >>
rect -5900 -20 -5800 0
rect -5900 -60 -5870 -20
rect -5830 -60 -5800 -20
rect -5900 -80 -5800 -60
rect -5700 -20 -5600 0
rect -5700 -60 -5670 -20
rect -5630 -60 -5600 -20
rect -5700 -80 -5600 -60
rect -4600 -20 -4500 0
rect -4600 -60 -4570 -20
rect -4530 -60 -4500 -20
rect -4600 -80 -4500 -60
rect -4400 -20 -4300 0
rect -4400 -60 -4370 -20
rect -4330 -60 -4300 -20
rect -4400 -80 -4300 -60
rect -3300 -20 -3200 0
rect -3300 -60 -3270 -20
rect -3230 -60 -3200 -20
rect -3300 -80 -3200 -60
rect -3100 -20 -3000 0
rect -3100 -60 -3070 -20
rect -3030 -60 -3000 -20
rect -3100 -80 -3000 -60
rect -2000 -20 -1900 0
rect -2000 -60 -1970 -20
rect -1930 -60 -1900 -20
rect -2000 -80 -1900 -60
rect -1800 -20 -1700 0
rect -1800 -60 -1770 -20
rect -1730 -60 -1700 -20
rect -1800 -80 -1700 -60
rect -700 -20 -600 0
rect -700 -60 -670 -20
rect -630 -60 -600 -20
rect -700 -80 -600 -60
rect -500 -20 -400 0
rect -500 -60 -470 -20
rect -430 -60 -400 -20
rect -500 -80 -400 -60
rect 100 -20 200 0
rect 100 -60 130 -20
rect 170 -60 200 -20
rect 100 -80 200 -60
rect 300 -20 400 0
rect 300 -60 330 -20
rect 370 -60 400 -20
rect 300 -80 400 -60
rect 1400 -20 1500 0
rect 1400 -60 1430 -20
rect 1470 -60 1500 -20
rect 1400 -80 1500 -60
rect 1600 -20 1700 0
rect 1600 -60 1630 -20
rect 1670 -60 1700 -20
rect 1600 -80 1700 -60
rect 2700 -20 2800 0
rect 2700 -60 2730 -20
rect 2770 -60 2800 -20
rect 2700 -80 2800 -60
rect 2900 -20 3000 0
rect 2900 -60 2930 -20
rect 2970 -60 3000 -20
rect 2900 -80 3000 -60
rect 4000 -20 4100 0
rect 4000 -60 4030 -20
rect 4070 -60 4100 -20
rect 4000 -80 4100 -60
rect 4200 -20 4300 0
rect 4200 -60 4230 -20
rect 4270 -60 4300 -20
rect 4200 -80 4300 -60
rect 5300 -20 5400 0
rect 5300 -60 5330 -20
rect 5370 -60 5400 -20
rect 5300 -80 5400 -60
rect 5500 -20 5600 0
rect 5500 -60 5530 -20
rect 5570 -60 5600 -20
rect 5500 -80 5600 -60
<< polycont >>
rect -5870 -60 -5830 -20
rect -5670 -60 -5630 -20
rect -4570 -60 -4530 -20
rect -4370 -60 -4330 -20
rect -3270 -60 -3230 -20
rect -3070 -60 -3030 -20
rect -1970 -60 -1930 -20
rect -1770 -60 -1730 -20
rect -670 -60 -630 -20
rect -470 -60 -430 -20
rect 130 -60 170 -20
rect 330 -60 370 -20
rect 1430 -60 1470 -20
rect 1630 -60 1670 -20
rect 2730 -60 2770 -20
rect 2930 -60 2970 -20
rect 4030 -60 4070 -20
rect 4230 -60 4270 -20
rect 5330 -60 5370 -20
rect 5530 -60 5570 -20
<< locali >>
rect -7160 2790 -7120 16450
rect -7080 5420 -7040 16450
rect -7000 8050 -6960 16450
rect -6920 10680 -6880 16450
rect -5040 16430 -4960 16450
rect -5040 16390 -5020 16430
rect -4980 16390 -4960 16430
rect -5040 16200 -4960 16390
rect -5040 16160 -5020 16200
rect -4980 16160 -4960 16200
rect -5040 16140 -4960 16160
rect -4180 15940 -4140 16450
rect -4100 16060 -4060 16450
rect -4020 16140 -3980 16450
rect -3940 16220 -3900 16450
rect -3740 16430 -3660 16450
rect -3740 16390 -3720 16430
rect -3680 16390 -3660 16430
rect -3940 16180 -3860 16220
rect -4020 16100 -3940 16140
rect -4100 16040 -4020 16060
rect -4100 16000 -4080 16040
rect -4040 16000 -4020 16040
rect -4100 15980 -4020 16000
rect -3980 16020 -3940 16100
rect -3900 16100 -3860 16180
rect -3740 16200 -3660 16390
rect -2440 16430 -2360 16450
rect -2440 16390 -2420 16430
rect -2380 16390 -2360 16430
rect -3740 16160 -3720 16200
rect -3680 16160 -3660 16200
rect -3740 16140 -3660 16160
rect -3120 16180 -2640 16220
rect -3120 16100 -3080 16180
rect -2800 16120 -2720 16140
rect -2800 16100 -2780 16120
rect -3900 16060 -3080 16100
rect -3040 16080 -2780 16100
rect -2740 16080 -2720 16120
rect -3040 16060 -2720 16080
rect -2680 16100 -2640 16180
rect -2440 16200 -2360 16390
rect -1140 16430 -1060 16450
rect -1140 16390 -1120 16430
rect -1080 16390 -1060 16430
rect -2440 16160 -2420 16200
rect -2380 16160 -2360 16200
rect -2440 16140 -2360 16160
rect -1820 16200 -1420 16220
rect -1820 16180 -1480 16200
rect -1820 16100 -1780 16180
rect -1500 16160 -1480 16180
rect -1440 16160 -1420 16200
rect -1500 16140 -1420 16160
rect -1140 16200 -1060 16390
rect -1140 16160 -1120 16200
rect -1080 16160 -1060 16200
rect -1140 16140 -1060 16160
rect 760 16430 840 16450
rect 760 16390 780 16430
rect 820 16390 840 16430
rect 760 16200 840 16390
rect 760 16160 780 16200
rect 820 16160 840 16200
rect 760 16140 840 16160
rect 2060 16430 2140 16450
rect 2060 16390 2080 16430
rect 2120 16390 2140 16430
rect 2060 16200 2140 16390
rect 2060 16160 2080 16200
rect 2120 16160 2140 16200
rect 2060 16140 2140 16160
rect 3360 16430 3440 16450
rect 3360 16390 3380 16430
rect 3420 16390 3440 16430
rect 3360 16200 3440 16390
rect 3360 16160 3380 16200
rect 3420 16160 3440 16200
rect 3360 16140 3440 16160
rect 4660 16430 4740 16450
rect 4660 16390 4680 16430
rect 4720 16390 4740 16430
rect 4660 16200 4740 16390
rect 4660 16160 4680 16200
rect 4720 16160 4740 16200
rect 4660 16140 4740 16160
rect 5960 16430 6040 16450
rect 5960 16390 5980 16430
rect 6020 16390 6040 16430
rect 5960 16200 6040 16390
rect 5960 16160 5980 16200
rect 6020 16160 6040 16200
rect 5960 16140 6040 16160
rect -2680 16060 -1780 16100
rect -1740 16060 280 16100
rect -3040 16020 -3000 16060
rect -1740 16020 -1700 16060
rect 240 16020 280 16060
rect -3980 15980 -3000 16020
rect -2960 15980 -1700 16020
rect -1660 15980 200 16020
rect 240 15980 1420 16020
rect -2960 15940 -2920 15980
rect -1660 15940 -1620 15980
rect 160 15940 200 15980
rect 1380 15940 1420 15980
rect -4180 15900 -2920 15940
rect -2880 15900 -1620 15940
rect -1580 15900 120 15940
rect 160 15900 1340 15940
rect 1380 15900 2640 15940
rect -4180 15860 -4140 15900
rect -2880 15860 -2840 15900
rect -1580 15860 -1540 15900
rect 80 15860 120 15900
rect 1300 15860 1340 15900
rect 2600 15860 2640 15900
rect -6840 15840 -6760 15860
rect -6840 15800 -6820 15840
rect -6780 15800 -6760 15840
rect -6840 15780 -6760 15800
rect -6700 15840 -6620 15860
rect -6700 15800 -6680 15840
rect -6640 15800 -6620 15840
rect -6700 15780 -6620 15800
rect -5400 15840 -4140 15860
rect -5400 15800 -5380 15840
rect -5340 15820 -4140 15840
rect -4100 15840 -2840 15860
rect -5340 15800 -5320 15820
rect -5400 15780 -5320 15800
rect -4100 15800 -4080 15840
rect -4040 15820 -2840 15840
rect -2800 15840 -1540 15860
rect -4040 15800 -4020 15820
rect -4100 15780 -4020 15800
rect -2800 15800 -2780 15840
rect -2740 15820 -1540 15840
rect -1500 15840 0 15860
rect -2740 15800 -2720 15820
rect -2800 15780 -2720 15800
rect -1500 15800 -1480 15840
rect -1440 15820 0 15840
rect 80 15820 1260 15860
rect 1300 15820 2560 15860
rect 2600 15820 3860 15860
rect -1440 15800 -1420 15820
rect -1500 15780 -1420 15800
rect -6840 13310 -6800 15780
rect -40 15700 0 15820
rect 1220 15780 1260 15820
rect 2520 15780 2560 15820
rect 3820 15780 3860 15820
rect -260 15620 0 15660
rect -260 13310 -220 15620
rect -6840 13270 -6760 13310
rect -300 13270 -220 13310
rect -120 13010 0 13030
rect -120 12970 -100 13010
rect -60 12990 0 13010
rect -60 12970 -40 12990
rect -120 12950 -40 12970
rect -6920 10640 -6760 10680
rect -300 10660 -190 10680
rect -300 10640 -250 10660
rect -270 10620 -250 10640
rect -210 10620 -190 10660
rect -270 10600 -190 10620
rect -270 10380 0 10400
rect -270 10340 -250 10380
rect -210 10360 0 10380
rect -210 10340 -190 10360
rect -270 10320 -190 10340
rect -7000 8010 -6760 8050
rect -300 8010 -220 8050
rect -260 7770 -220 8010
rect -260 7730 0 7770
rect -270 5440 -190 5460
rect -270 5420 -250 5440
rect -7080 5380 -6760 5420
rect -300 5400 -250 5420
rect -210 5400 -190 5440
rect -300 5380 -190 5400
rect -190 5160 -110 5180
rect -190 5120 -170 5160
rect -130 5140 -110 5160
rect -130 5120 0 5140
rect -190 5100 0 5120
rect -130 2810 -50 2830
rect -130 2790 -110 2810
rect -7160 2750 -6760 2790
rect -300 2770 -110 2790
rect -70 2770 -50 2810
rect -300 2750 -50 2770
rect -260 2470 0 2510
rect -260 160 -220 2470
rect -6940 140 -6760 160
rect -6940 100 -6920 140
rect -6880 120 -6760 140
rect -300 120 -220 160
rect -6880 100 -6860 120
rect -6940 80 -6860 100
rect -6560 -20 -6480 0
rect -6560 -60 -6540 -20
rect -6500 -60 -6480 -20
rect -6560 -280 -6480 -60
rect -6560 -320 -6540 -280
rect -6500 -320 -6480 -280
rect -6560 -340 -6480 -320
rect -5890 -20 -5810 0
rect -5890 -60 -5870 -20
rect -5830 -60 -5810 -20
rect -5890 -520 -5810 -60
rect -5690 -20 -5610 0
rect -5690 -60 -5670 -20
rect -5630 -60 -5610 -20
rect -5690 -400 -5610 -60
rect -5260 -20 -5180 0
rect -5260 -60 -5240 -20
rect -5200 -60 -5180 -20
rect -5260 -280 -5180 -60
rect -5260 -320 -5240 -280
rect -5200 -320 -5180 -280
rect -5260 -340 -5180 -320
rect -4590 -20 -4510 0
rect -4590 -60 -4570 -20
rect -4530 -60 -4510 -20
rect -5690 -440 -5670 -400
rect -5630 -440 -5610 -400
rect -5690 -460 -5610 -440
rect -5890 -560 -5870 -520
rect -5830 -560 -5810 -520
rect -5890 -580 -5810 -560
rect -4590 -520 -4510 -60
rect -4390 -20 -4310 0
rect -4390 -60 -4370 -20
rect -4330 -60 -4310 -20
rect -4390 -400 -4310 -60
rect -3960 -20 -3880 0
rect -3960 -60 -3940 -20
rect -3900 -60 -3880 -20
rect -3960 -280 -3880 -60
rect -3960 -320 -3940 -280
rect -3900 -320 -3880 -280
rect -3960 -340 -3880 -320
rect -3290 -20 -3210 0
rect -3290 -60 -3270 -20
rect -3230 -60 -3210 -20
rect -4390 -440 -4370 -400
rect -4330 -440 -4310 -400
rect -4390 -460 -4310 -440
rect -4590 -560 -4570 -520
rect -4530 -560 -4510 -520
rect -4590 -580 -4510 -560
rect -3290 -520 -3210 -60
rect -3090 -20 -3010 0
rect -3090 -60 -3070 -20
rect -3030 -60 -3010 -20
rect -3090 -400 -3010 -60
rect -2660 -20 -2580 0
rect -2660 -60 -2640 -20
rect -2600 -60 -2580 -20
rect -2660 -280 -2580 -60
rect -2660 -320 -2640 -280
rect -2600 -320 -2580 -280
rect -2660 -340 -2580 -320
rect -1990 -20 -1910 0
rect -1990 -60 -1970 -20
rect -1930 -60 -1910 -20
rect -3090 -440 -3070 -400
rect -3030 -440 -3010 -400
rect -3090 -460 -3010 -440
rect -3290 -560 -3270 -520
rect -3230 -560 -3210 -520
rect -3290 -580 -3210 -560
rect -1990 -520 -1910 -60
rect -1790 -20 -1710 0
rect -1790 -60 -1770 -20
rect -1730 -60 -1710 -20
rect -1790 -400 -1710 -60
rect -1360 -20 -1280 0
rect -1360 -60 -1340 -20
rect -1300 -60 -1280 -20
rect -1360 -280 -1280 -60
rect -1360 -320 -1340 -280
rect -1300 -320 -1280 -280
rect -1360 -340 -1280 -320
rect -690 -20 -610 0
rect -690 -60 -670 -20
rect -630 -60 -610 -20
rect -1790 -440 -1770 -400
rect -1730 -440 -1710 -400
rect -1790 -460 -1710 -440
rect -1990 -560 -1970 -520
rect -1930 -560 -1910 -520
rect -1990 -580 -1910 -560
rect -690 -520 -610 -60
rect -490 -20 -410 0
rect -490 -60 -470 -20
rect -430 -60 -410 -20
rect -490 -400 -410 -60
rect -490 -440 -470 -400
rect -430 -440 -410 -400
rect -490 -460 -410 -440
rect 110 -20 190 0
rect 110 -60 130 -20
rect 170 -60 190 -20
rect 110 -400 190 -60
rect 110 -440 130 -400
rect 170 -440 190 -400
rect 110 -460 190 -440
rect 310 -20 390 0
rect 310 -60 330 -20
rect 370 -60 390 -20
rect -690 -560 -670 -520
rect -630 -560 -610 -520
rect -690 -580 -610 -560
rect 310 -520 390 -60
rect 1010 -20 1090 0
rect 1010 -60 1030 -20
rect 1070 -60 1090 -20
rect 1010 -280 1090 -60
rect 1010 -320 1030 -280
rect 1070 -320 1090 -280
rect 1010 -340 1090 -320
rect 1410 -20 1490 0
rect 1410 -60 1430 -20
rect 1470 -60 1490 -20
rect 1410 -400 1490 -60
rect 1410 -440 1430 -400
rect 1470 -440 1490 -400
rect 1410 -460 1490 -440
rect 1610 -20 1690 0
rect 1610 -60 1630 -20
rect 1670 -60 1690 -20
rect 310 -560 330 -520
rect 370 -560 390 -520
rect 310 -580 390 -560
rect 1610 -520 1690 -60
rect 2310 -20 2390 0
rect 2310 -60 2330 -20
rect 2370 -60 2390 -20
rect 2310 -280 2390 -60
rect 2310 -320 2330 -280
rect 2370 -320 2390 -280
rect 2310 -340 2390 -320
rect 2710 -20 2790 0
rect 2710 -60 2730 -20
rect 2770 -60 2790 -20
rect 2710 -400 2790 -60
rect 2710 -440 2730 -400
rect 2770 -440 2790 -400
rect 2710 -460 2790 -440
rect 2910 -20 2990 0
rect 2910 -60 2930 -20
rect 2970 -60 2990 -20
rect 1610 -560 1630 -520
rect 1670 -560 1690 -520
rect 1610 -580 1690 -560
rect 2910 -520 2990 -60
rect 3610 -20 3690 0
rect 3610 -60 3630 -20
rect 3670 -60 3690 -20
rect 3610 -280 3690 -60
rect 3610 -320 3630 -280
rect 3670 -320 3690 -280
rect 3610 -340 3690 -320
rect 4010 -20 4090 0
rect 4010 -60 4030 -20
rect 4070 -60 4090 -20
rect 4010 -400 4090 -60
rect 4010 -440 4030 -400
rect 4070 -440 4090 -400
rect 4010 -460 4090 -440
rect 4210 -20 4290 0
rect 4210 -60 4230 -20
rect 4270 -60 4290 -20
rect 2910 -560 2930 -520
rect 2970 -560 2990 -520
rect 2910 -580 2990 -560
rect 4210 -520 4290 -60
rect 4910 -20 4990 0
rect 4910 -60 4930 -20
rect 4970 -60 4990 -20
rect 4910 -280 4990 -60
rect 4910 -320 4930 -280
rect 4970 -320 4990 -280
rect 4910 -340 4990 -320
rect 5310 -20 5390 0
rect 5310 -60 5330 -20
rect 5370 -60 5390 -20
rect 5310 -400 5390 -60
rect 5310 -440 5330 -400
rect 5370 -440 5390 -400
rect 5310 -460 5390 -440
rect 5510 -20 5590 0
rect 5510 -60 5530 -20
rect 5570 -60 5590 -20
rect 4210 -560 4230 -520
rect 4270 -560 4290 -520
rect 4210 -580 4290 -560
rect 5510 -520 5590 -60
rect 6210 -20 6290 0
rect 6210 -60 6230 -20
rect 6270 -60 6290 -20
rect 6210 -280 6290 -60
rect 6210 -320 6230 -280
rect 6270 -320 6290 -280
rect 6210 -340 6290 -320
rect 5510 -560 5530 -520
rect 5570 -560 5590 -520
rect 5510 -580 5590 -560
<< viali >>
rect -5020 16390 -4980 16430
rect -5020 16160 -4980 16200
rect -3720 16390 -3680 16430
rect -4080 16000 -4040 16040
rect -2420 16390 -2380 16430
rect -3720 16160 -3680 16200
rect -2780 16080 -2740 16120
rect -1120 16390 -1080 16430
rect -2420 16160 -2380 16200
rect -1480 16160 -1440 16200
rect -1120 16160 -1080 16200
rect 780 16390 820 16430
rect 780 16160 820 16200
rect 2080 16390 2120 16430
rect 2080 16160 2120 16200
rect 3380 16390 3420 16430
rect 3380 16160 3420 16200
rect 4680 16390 4720 16430
rect 4680 16160 4720 16200
rect 5980 16390 6020 16430
rect 5980 16160 6020 16200
rect -6820 15800 -6780 15840
rect -6680 15800 -6640 15840
rect -5380 15800 -5340 15840
rect -4080 15800 -4040 15840
rect -2780 15800 -2740 15840
rect -1480 15800 -1440 15840
rect -100 12970 -60 13010
rect -250 10620 -210 10660
rect -250 10340 -210 10380
rect -250 5400 -210 5440
rect -170 5120 -130 5160
rect -110 2770 -70 2810
rect -6920 100 -6880 140
rect -6540 -60 -6500 -20
rect -6540 -320 -6500 -280
rect -5240 -60 -5200 -20
rect -5240 -320 -5200 -280
rect -5670 -440 -5630 -400
rect -5870 -560 -5830 -520
rect -3940 -60 -3900 -20
rect -3940 -320 -3900 -280
rect -4370 -440 -4330 -400
rect -4570 -560 -4530 -520
rect -2640 -60 -2600 -20
rect -2640 -320 -2600 -280
rect -3070 -440 -3030 -400
rect -3270 -560 -3230 -520
rect -1340 -60 -1300 -20
rect -1340 -320 -1300 -280
rect -1770 -440 -1730 -400
rect -1970 -560 -1930 -520
rect -470 -440 -430 -400
rect 130 -440 170 -400
rect -670 -560 -630 -520
rect 1030 -60 1070 -20
rect 1030 -320 1070 -280
rect 1430 -440 1470 -400
rect 330 -560 370 -520
rect 2330 -60 2370 -20
rect 2330 -320 2370 -280
rect 2730 -440 2770 -400
rect 1630 -560 1670 -520
rect 3630 -60 3670 -20
rect 3630 -320 3670 -280
rect 4030 -440 4070 -400
rect 2930 -560 2970 -520
rect 4930 -60 4970 -20
rect 4930 -320 4970 -280
rect 5330 -440 5370 -400
rect 4230 -560 4270 -520
rect 6230 -60 6270 -20
rect 6230 -320 6270 -280
rect 5530 -560 5570 -520
<< metal1 >>
rect -7300 -520 -7240 16450
rect -7180 -400 -7120 16450
rect -7060 -260 -7000 16450
rect -6920 15860 -6860 16450
rect -5040 16430 -4960 16450
rect -3740 16430 -3660 16450
rect -2440 16430 -2360 16450
rect -1140 16430 -1060 16450
rect 760 16430 840 16450
rect 2060 16430 2140 16450
rect 3360 16430 3440 16450
rect 4660 16430 4740 16450
rect 5960 16430 6040 16450
rect -6330 16390 -5020 16430
rect -4980 16390 -3720 16430
rect -3680 16390 -2420 16430
rect -2380 16390 -1120 16430
rect -1080 16390 780 16430
rect 820 16390 2080 16430
rect 2120 16390 3380 16430
rect 3420 16390 4680 16430
rect 4720 16390 5980 16430
rect 6020 16390 6560 16430
rect -6330 16370 6560 16390
rect -6920 15840 -6620 15860
rect -6920 15800 -6820 15840
rect -6780 15800 -6680 15840
rect -6640 15800 -6620 15840
rect -6920 15780 -6620 15800
rect -6330 15780 -6270 16370
rect -5900 16250 6560 16310
rect -5900 15780 -5840 16250
rect -5040 16200 -4960 16220
rect -5040 16160 -5020 16200
rect -4980 16160 -4960 16200
rect -5040 16140 -4960 16160
rect -5400 15840 -5320 15860
rect -5400 15800 -5380 15840
rect -5340 15800 -5320 15840
rect -5400 15780 -5320 15800
rect -5030 15780 -4970 16140
rect -4600 15780 -4540 16250
rect -3740 16200 -3660 16220
rect -3740 16160 -3720 16200
rect -3680 16160 -3660 16200
rect -3740 16140 -3660 16160
rect -4100 16040 -4020 16060
rect -4100 16000 -4080 16040
rect -4040 16000 -4020 16040
rect -4100 15980 -4020 16000
rect -4050 15860 -4020 15980
rect -4100 15840 -4020 15860
rect -4100 15800 -4080 15840
rect -4040 15800 -4020 15840
rect -4100 15780 -4020 15800
rect -3730 15780 -3670 16140
rect -3300 15780 -3240 16250
rect -2440 16200 -2360 16220
rect -2440 16160 -2420 16200
rect -2380 16160 -2360 16200
rect -2440 16140 -2360 16160
rect -2800 16120 -2720 16140
rect -2800 16080 -2780 16120
rect -2740 16080 -2720 16120
rect -2800 16060 -2720 16080
rect -2750 15860 -2720 16060
rect -2800 15840 -2720 15860
rect -2800 15800 -2780 15840
rect -2740 15800 -2720 15840
rect -2800 15780 -2720 15800
rect -2430 15780 -2370 16140
rect -2000 15780 -1940 16250
rect -1500 16200 -1420 16220
rect -1500 16160 -1480 16200
rect -1440 16160 -1420 16200
rect -1500 16140 -1420 16160
rect -1140 16200 -1060 16220
rect -1140 16160 -1120 16200
rect -1080 16160 -1060 16200
rect -1140 16140 -1060 16160
rect -1450 15860 -1420 16140
rect -1500 15840 -1420 15860
rect -1500 15800 -1480 15840
rect -1440 15800 -1420 15840
rect -1500 15780 -1420 15800
rect -1130 15780 -1070 16140
rect -700 15780 -640 16250
rect 340 15780 400 16250
rect 760 16200 840 16220
rect 760 16160 780 16200
rect 820 16160 840 16200
rect 760 16140 840 16160
rect 770 15780 830 16140
rect 1640 15780 1700 16250
rect 2060 16200 2140 16220
rect 2060 16160 2080 16200
rect 2120 16160 2140 16200
rect 2060 16140 2140 16160
rect 2070 15780 2130 16140
rect 2940 15780 3000 16250
rect 3360 16200 3440 16220
rect 3360 16160 3380 16200
rect 3420 16160 3440 16200
rect 3360 16140 3440 16160
rect 3370 15780 3430 16140
rect 4240 15780 4300 16250
rect 4660 16200 4740 16220
rect 4660 16160 4680 16200
rect 4720 16160 4740 16200
rect 4660 16140 4740 16160
rect 4670 15780 4730 16140
rect 5540 15780 5600 16250
rect 5960 16200 6040 16220
rect 5960 16160 5980 16200
rect 6020 16160 6040 16200
rect 5960 16140 6040 16160
rect 5970 15780 6030 16140
rect -6920 13230 -6860 15780
rect -6920 13150 -6800 13230
rect -6920 10600 -6860 13150
rect -120 13010 -40 13030
rect -120 12970 -100 13010
rect -60 12970 -40 13010
rect -120 12950 -40 12970
rect -270 10660 -190 10680
rect -270 10620 -250 10660
rect -210 10630 -190 10660
rect -210 10620 -130 10630
rect -270 10600 -130 10620
rect -6920 10520 -6800 10600
rect -6920 7970 -6860 10520
rect -270 10380 -190 10400
rect -270 10340 -250 10380
rect -210 10340 -190 10380
rect -270 10320 -190 10340
rect -6920 7890 -6800 7970
rect -6920 5340 -6860 7890
rect -270 5460 -240 10320
rect -270 5440 -190 5460
rect -270 5400 -250 5440
rect -210 5400 -190 5440
rect -270 5380 -190 5400
rect -6920 5260 -6800 5340
rect -6920 2710 -6860 5260
rect -160 5180 -130 10600
rect -190 5160 -110 5180
rect -190 5120 -170 5160
rect -130 5120 -110 5160
rect -190 5100 -110 5120
rect -80 2830 -50 12950
rect -130 2810 -50 2830
rect -130 2770 -110 2810
rect -70 2770 -50 2810
rect -130 2750 -50 2770
rect -6920 2630 -6800 2710
rect -6920 160 -6860 2630
rect -6940 140 -6860 160
rect -6940 100 -6920 140
rect -6880 100 -6860 140
rect -6940 80 -6860 100
rect -6920 0 -6800 80
rect -6920 -140 -6860 0
rect -6570 -20 -6480 0
rect -6570 -60 -6540 -20
rect -6500 -60 -6480 -20
rect -6560 -80 -6480 -60
rect -6450 -140 -6390 0
rect -5590 -140 -5530 0
rect -5270 -20 -5180 0
rect -5270 -60 -5240 -20
rect -5200 -60 -5180 -20
rect -5260 -80 -5180 -60
rect -5150 -140 -5090 0
rect -4290 -140 -4230 0
rect -3970 -20 -3880 0
rect -3970 -60 -3940 -20
rect -3900 -60 -3880 -20
rect -3960 -80 -3880 -60
rect -3850 -140 -3790 0
rect -2990 -140 -2930 0
rect -2670 -20 -2580 0
rect -2670 -60 -2640 -20
rect -2600 -60 -2580 -20
rect -2660 -80 -2580 -60
rect -2550 -140 -2490 0
rect -1690 -140 -1630 0
rect -1370 -20 -1280 0
rect -1370 -60 -1340 -20
rect -1300 -60 -1280 -20
rect -1360 -80 -1280 -60
rect -1250 -140 -1190 0
rect -390 -140 -330 0
rect 30 -140 90 0
rect 890 -140 950 0
rect 1010 -20 1090 0
rect 1010 -60 1030 -20
rect 1070 -60 1090 -20
rect 1010 -80 1090 -60
rect 1330 -140 1390 0
rect 2190 -140 2250 0
rect 2310 -20 2390 0
rect 2310 -60 2330 -20
rect 2370 -60 2390 -20
rect 2310 -80 2390 -60
rect 2630 -140 2690 0
rect 3490 -140 3550 0
rect 3610 -20 3690 0
rect 3610 -60 3630 -20
rect 3670 -60 3690 -20
rect 3610 -80 3690 -60
rect 3930 -140 3990 0
rect 4790 -140 4850 0
rect 4910 -20 4990 0
rect 4910 -60 4930 -20
rect 4970 -60 4990 -20
rect 4910 -80 4990 -60
rect 5230 -140 5290 0
rect 6090 -140 6150 0
rect 6210 -20 6290 0
rect 6210 -60 6230 -20
rect 6270 -60 6290 -20
rect 6210 -80 6290 -60
rect 6320 -140 6350 0
rect 6500 -140 6560 15780
rect -6920 -200 6560 -140
rect -7060 -280 6560 -260
rect -7060 -320 -6540 -280
rect -6500 -320 -5240 -280
rect -5200 -320 -3940 -280
rect -3900 -320 -2640 -280
rect -2600 -320 -1340 -280
rect -1300 -320 1030 -280
rect 1070 -320 2330 -280
rect 2370 -320 3630 -280
rect 3670 -320 4930 -280
rect 4970 -320 6230 -280
rect 6270 -320 6560 -280
rect -6560 -340 -6480 -320
rect -5260 -340 -5180 -320
rect -3960 -340 -3880 -320
rect -2660 -340 -2580 -320
rect -1360 -340 -1280 -320
rect 1010 -340 1090 -320
rect 2310 -340 2390 -320
rect 3610 -340 3690 -320
rect 4910 -340 4990 -320
rect 6210 -340 6290 -320
rect -5690 -400 -5610 -380
rect -4390 -400 -4310 -380
rect -3090 -400 -3010 -380
rect -1790 -400 -1710 -380
rect -490 -400 -410 -380
rect 110 -400 190 -380
rect 1410 -400 1490 -380
rect 2710 -400 2790 -380
rect 4010 -400 4090 -380
rect 5310 -400 5390 -380
rect -7180 -440 -5670 -400
rect -5630 -440 -4370 -400
rect -4330 -440 -3070 -400
rect -3030 -440 -1770 -400
rect -1730 -440 -470 -400
rect -430 -440 130 -400
rect 170 -440 1430 -400
rect 1470 -440 2730 -400
rect 2770 -440 4030 -400
rect 4070 -440 5330 -400
rect 5370 -440 6560 -400
rect -7180 -460 6560 -440
rect -5890 -520 -5810 -500
rect -4590 -520 -4510 -500
rect -3290 -520 -3210 -500
rect -1990 -520 -1910 -500
rect -690 -520 -610 -500
rect 310 -520 390 -500
rect 1610 -520 1690 -500
rect 2910 -520 2990 -500
rect 4210 -520 4290 -500
rect 5510 -520 5590 -500
rect -7300 -560 -5870 -520
rect -5830 -560 -4570 -520
rect -4530 -560 -3270 -520
rect -3230 -560 -1970 -520
rect -1930 -560 -670 -520
rect -630 -560 330 -520
rect 370 -560 1630 -520
rect 1670 -560 2930 -520
rect 2970 -560 4230 -520
rect 4270 -560 5530 -520
rect 5570 -560 6560 -520
rect -7300 -580 6560 -560
use half_dac_for_mirroring  half_dac_for_mirroring_0
timestamp 1702591987
transform 1 0 1300 0 1 2630
box -1396 -2630 5325 13211
use half_dac_for_mirroring  half_dac_for_mirroring_1
timestamp 1702591987
transform -1 0 -1600 0 -1 13150
box -1396 -2630 5325 13211
<< labels >>
flabel locali -3920 16450 -3920 16450 1 FreeSans 320 0 0 0 X0
port 1 n
flabel locali -4000 16450 -4000 16450 1 FreeSans 320 0 0 0 X1
port 2 n
flabel locali -4080 16450 -4080 16450 1 FreeSans 320 0 0 0 X2
port 3 n
flabel locali -4160 16450 -4160 16450 1 FreeSans 320 0 0 0 X3
port 4 n
flabel locali -6900 16450 -6900 16450 1 FreeSans 320 0 0 0 Y0
port 5 n
flabel locali -6980 16450 -6980 16450 1 FreeSans 320 0 0 0 Y1
port 6 n
flabel locali -7060 16450 -7060 16450 1 FreeSans 320 0 0 0 Y2
port 7 n
flabel locali -7140 16450 -7140 16450 1 FreeSans 320 0 0 0 Y3
port 8 n
flabel metal1 6560 16280 6560 16280 3 FreeSans 320 0 0 0 I1
port 9 e
flabel metal1 6560 16400 6560 16400 3 FreeSans 320 0 0 0 I2
port 10 e
flabel metal1 6560 -290 6560 -290 3 FreeSans 320 0 0 0 VDD
port 11 e
flabel metal1 6560 -170 6560 -170 3 FreeSans 320 0 0 0 GND
port 12 e
flabel metal1 6560 -430 6560 -430 3 FreeSans 480 0 0 0 Vbn
port 13 e
flabel metal1 6560 -550 6560 -550 3 FreeSans 480 0 0 0 Vcn
port 14 e
<< end >>
