magic
tech sky130A
timestamp 1702266255
<< nwell >>
rect 430 765 570 1245
<< nmos >>
rect 50 0 100 1200
rect 150 0 200 1200
rect 280 1160 380 1175
rect 280 1095 380 1110
rect 280 1030 380 1045
rect 280 835 380 850
rect 260 405 310 705
rect 260 0 310 300
<< pmos >>
rect 450 1160 550 1175
rect 450 1095 550 1110
rect 450 1030 550 1045
rect 450 835 550 850
<< ndiff >>
rect 0 0 50 1200
rect 100 0 150 1200
rect 200 705 250 1200
rect 280 1175 380 1225
rect 280 1110 380 1160
rect 280 1045 380 1095
rect 280 980 380 1030
rect 280 850 380 900
rect 280 785 380 835
rect 200 405 260 705
rect 310 405 360 705
rect 200 300 250 405
rect 200 0 260 300
rect 310 0 360 300
<< pdiff >>
rect 450 1175 550 1225
rect 450 1110 550 1160
rect 450 1045 550 1095
rect 450 980 550 1030
rect 450 850 550 900
rect 450 785 550 835
<< psubdiff >>
rect 280 935 380 950
rect 280 915 295 935
rect 365 915 380 935
rect 280 900 380 915
<< nsubdiff >>
rect 450 935 550 950
rect 450 915 465 935
rect 535 915 550 935
rect 450 900 550 915
<< psubdiffcont >>
rect 295 915 365 935
<< nsubdiffcont >>
rect 465 915 535 935
<< poly >>
rect 50 1200 100 1215
rect 150 1200 200 1215
rect 395 1175 435 1195
rect 265 1160 280 1175
rect 380 1160 450 1175
rect 550 1160 565 1175
rect 395 1155 435 1160
rect 395 1110 435 1130
rect 265 1095 280 1110
rect 380 1095 450 1110
rect 550 1095 565 1110
rect 395 1090 435 1095
rect 395 1045 435 1065
rect 265 1030 280 1045
rect 380 1030 450 1045
rect 550 1030 565 1045
rect 395 1025 435 1030
rect 395 865 435 875
rect 395 850 405 865
rect 265 835 280 850
rect 380 845 405 850
rect 425 850 435 865
rect 425 845 450 850
rect 380 835 450 845
rect 550 835 565 850
rect 260 755 310 770
rect 260 735 275 755
rect 295 735 310 755
rect 260 705 310 735
rect 260 390 310 405
rect 260 350 310 365
rect 260 330 275 350
rect 295 330 310 350
rect 260 300 310 330
rect 50 -15 100 0
rect 150 -15 200 0
rect 260 -15 310 0
<< polycont >>
rect 405 845 425 865
rect 275 735 295 755
rect 275 330 295 350
<< locali >>
rect 285 1200 375 1220
rect 245 1180 375 1200
rect 455 1200 545 1220
rect 245 1025 265 1180
rect 395 1155 435 1195
rect 455 1180 585 1200
rect 455 1145 545 1155
rect 395 1090 435 1130
rect 455 1125 465 1145
rect 535 1125 545 1145
rect 455 1115 545 1125
rect 565 1090 585 1180
rect 285 1080 375 1090
rect 285 1060 295 1080
rect 365 1060 375 1080
rect 455 1070 585 1090
rect 285 1050 375 1060
rect 395 1025 435 1065
rect 455 1050 545 1070
rect 245 1005 375 1025
rect 455 1005 545 1025
rect 245 765 265 1005
rect 285 985 545 1005
rect 285 935 375 945
rect 285 915 295 935
rect 365 915 375 935
rect 285 885 375 915
rect 285 865 295 885
rect 365 865 375 885
rect 405 875 425 985
rect 455 935 545 945
rect 455 915 465 935
rect 535 915 545 935
rect 455 885 545 915
rect 285 855 375 865
rect 395 865 435 875
rect 395 845 405 865
rect 425 845 435 865
rect 455 865 465 885
rect 535 865 545 885
rect 455 855 545 865
rect 395 835 435 845
rect 285 810 375 830
rect 455 810 545 830
rect 285 790 545 810
rect 245 755 305 765
rect 245 745 275 755
rect 265 735 275 745
rect 295 735 305 755
rect 265 725 305 735
rect 315 690 355 700
rect 315 420 325 690
rect 345 420 355 690
rect 315 410 355 420
rect 375 360 395 790
rect 265 350 395 360
rect 265 330 275 350
rect 295 340 395 350
rect 295 330 305 340
rect 265 320 305 330
rect 315 285 355 295
rect 315 15 325 285
rect 345 15 355 285
rect 315 5 355 15
<< viali >>
rect 465 1125 535 1145
rect 295 1060 365 1080
rect 295 915 365 935
rect 295 865 365 885
rect 465 915 535 935
rect 465 865 535 885
rect 325 420 345 690
rect 325 15 345 285
<< metal1 >>
rect 455 1145 545 1155
rect 455 1125 465 1145
rect 535 1125 545 1145
rect 455 1115 545 1125
rect 285 1080 375 1090
rect 285 1060 295 1080
rect 365 1060 375 1080
rect 285 1050 375 1060
rect 285 935 375 945
rect 285 915 295 935
rect 365 915 375 935
rect 285 885 375 915
rect 285 865 295 885
rect 365 865 375 885
rect 285 855 375 865
rect 455 935 545 945
rect 455 915 465 935
rect 535 915 545 935
rect 455 885 545 915
rect 455 865 465 885
rect 535 865 545 885
rect 455 855 545 865
rect 315 690 355 700
rect 315 420 325 690
rect 345 420 355 690
rect 315 410 355 420
rect 315 285 355 295
rect 315 15 325 285
rect 345 15 355 285
rect 315 5 355 15
<< end >>
