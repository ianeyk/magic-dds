magic
tech sky130A
magscale 1 2
timestamp 1702743177
<< error_s >>
rect 4085 430 4100 630
rect 4110 430 4154 630
<< nwell >>
rect 500 620 510 630
rect 970 620 980 630
rect 1560 620 1580 630
rect 2170 620 2180 630
rect 2890 620 2910 630
rect 3490 620 3510 630
rect 490 440 530 620
rect 960 440 1000 620
rect 1560 440 1600 620
rect 2160 440 2200 620
rect 2890 440 2930 620
rect 3490 440 3530 620
rect 500 430 510 440
rect 970 430 980 440
rect 1560 430 1580 440
rect 2170 430 2180 440
rect 2890 430 2910 440
rect 3490 430 3510 440
<< pdiff >>
rect 500 620 510 630
rect 970 620 980 630
rect 490 440 510 620
rect 960 440 980 620
rect 500 430 510 440
rect 970 430 980 440
rect 1560 430 1580 630
rect 2170 620 2180 630
rect 2160 440 2180 620
rect 2170 430 2180 440
rect 2890 430 2910 630
rect 3490 430 3510 630
<< nsubdiff >>
rect 510 440 530 620
rect 980 440 1000 620
rect 1580 440 1600 620
rect 2180 440 2200 620
rect 2910 440 2930 620
rect 3510 440 3530 620
<< poly >>
rect 240 -20 320 0
rect 240 -60 260 -20
rect 300 -60 320 -20
rect 240 -80 320 -60
rect 370 -280 400 0
rect 760 -200 790 0
rect 840 -80 870 0
rect 1230 -80 1260 10
rect 840 -100 920 -80
rect 840 -140 860 -100
rect 900 -140 920 -100
rect 840 -160 920 -140
rect 1180 -100 1260 -80
rect 1180 -140 1200 -100
rect 1240 -140 1260 -100
rect 1180 -160 1260 -140
rect 710 -220 790 -200
rect 710 -260 730 -220
rect 770 -260 790 -220
rect 710 -280 790 -260
rect 370 -300 450 -280
rect 370 -340 390 -300
rect 430 -340 450 -300
rect 370 -360 450 -340
rect 1310 -400 1340 0
rect 1260 -420 1340 -400
rect 1260 -460 1280 -420
rect 1320 -460 1340 -420
rect 1260 -480 1340 -460
rect 1390 -600 1420 0
rect 1830 -200 1860 10
rect 1780 -220 1860 -200
rect 1780 -260 1800 -220
rect 1840 -260 1860 -220
rect 1780 -280 1860 -260
rect 1910 -480 1940 0
rect 1860 -500 1940 -480
rect 1860 -540 1880 -500
rect 1920 -540 1940 -500
rect 1860 -560 1940 -540
rect 1390 -620 1470 -600
rect 1390 -660 1410 -620
rect 1450 -660 1470 -620
rect 1390 -680 1470 -660
rect 1990 -680 2020 0
rect 2430 -80 2460 0
rect 2380 -100 2460 -80
rect 2380 -140 2400 -100
rect 2440 -140 2460 -100
rect 2380 -160 2460 -140
rect 2510 -680 2540 0
rect 1970 -700 2050 -680
rect 1970 -740 1990 -700
rect 2030 -740 2050 -700
rect 1970 -760 2050 -740
rect 2460 -700 2540 -680
rect 2460 -740 2480 -700
rect 2520 -740 2540 -700
rect 2460 -760 2540 -740
rect 2590 -880 2620 0
rect 2530 -900 2620 -880
rect 2530 -940 2550 -900
rect 2590 -940 2620 -900
rect 2530 -960 2620 -940
rect 2670 -1080 2700 0
rect 3110 -20 3190 0
rect 3110 -60 3130 -20
rect 3170 -60 3190 -20
rect 3110 -80 3190 -60
rect 3240 -480 3270 30
rect 3190 -500 3270 -480
rect 3190 -540 3210 -500
rect 3250 -540 3270 -500
rect 3190 -560 3270 -540
rect 3320 -600 3350 0
rect 3760 -80 3790 0
rect 3710 -100 3790 -80
rect 3710 -140 3730 -100
rect 3770 -140 3790 -100
rect 3710 -150 3790 -140
rect 3840 -200 3870 60
rect 3790 -220 3870 -200
rect 3790 -260 3810 -220
rect 3850 -260 3870 -220
rect 3790 -280 3870 -260
rect 3320 -620 3400 -600
rect 3320 -660 3340 -620
rect 3380 -660 3400 -620
rect 3320 -680 3400 -660
rect 3920 -800 3950 0
rect 3920 -820 4000 -800
rect 3920 -860 3940 -820
rect 3980 -860 4000 -820
rect 3920 -880 4000 -860
rect 2600 -1100 2700 -1080
rect 2600 -1140 2620 -1100
rect 2660 -1140 2700 -1100
rect 2600 -1160 2700 -1140
<< polycont >>
rect 260 -60 300 -20
rect 860 -140 900 -100
rect 1200 -140 1240 -100
rect 730 -260 770 -220
rect 390 -340 430 -300
rect 1280 -460 1320 -420
rect 1800 -260 1840 -220
rect 1880 -540 1920 -500
rect 1410 -660 1450 -620
rect 2400 -140 2440 -100
rect 1990 -740 2030 -700
rect 2480 -740 2520 -700
rect 2550 -940 2590 -900
rect 3130 -60 3170 -20
rect 3210 -540 3250 -500
rect 3730 -140 3770 -100
rect 3810 -260 3850 -220
rect 3340 -660 3380 -620
rect 3940 -860 3980 -820
rect 2620 -1140 2660 -1100
<< locali >>
rect 490 440 530 620
rect 960 440 1000 620
rect 1560 440 1600 620
rect 2160 440 2200 620
rect 2890 440 2930 620
rect 3490 440 3530 620
rect 0 -20 7880 0
rect 0 -40 260 -20
rect 240 -60 260 -40
rect 300 -40 3130 -20
rect 300 -60 320 -40
rect 240 -80 320 -60
rect 3110 -60 3130 -40
rect 3170 -40 7880 -20
rect 3170 -60 3190 -40
rect 3110 -80 3190 -60
rect 840 -100 920 -80
rect 840 -120 860 -100
rect 0 -140 860 -120
rect 900 -120 920 -100
rect 1180 -100 1260 -80
rect 1180 -120 1200 -100
rect 900 -140 1200 -120
rect 1240 -120 1260 -100
rect 2380 -100 2460 -80
rect 2380 -120 2400 -100
rect 1240 -140 2400 -120
rect 2440 -120 2460 -100
rect 3710 -100 3790 -80
rect 3710 -120 3730 -100
rect 2440 -140 3730 -120
rect 3770 -120 3790 -100
rect 3770 -140 7880 -120
rect 0 -160 7880 -140
rect 0 -220 7880 -200
rect 0 -240 730 -220
rect 710 -260 730 -240
rect 770 -240 1800 -220
rect 770 -260 790 -240
rect 710 -280 790 -260
rect 1780 -260 1800 -240
rect 1840 -240 3810 -220
rect 1840 -260 1860 -240
rect 1780 -280 1860 -260
rect 3790 -260 3810 -240
rect 3850 -240 7880 -220
rect 3850 -260 3870 -240
rect 3790 -280 3870 -260
rect 370 -300 450 -280
rect 370 -320 390 -300
rect 0 -340 390 -320
rect 430 -320 450 -300
rect 430 -340 7880 -320
rect 0 -360 7880 -340
rect 0 -420 7880 -400
rect 0 -440 1280 -420
rect 1260 -460 1280 -440
rect 1320 -440 7880 -420
rect 1320 -460 1340 -440
rect 1260 -480 1340 -460
rect 1860 -500 1940 -480
rect 1860 -520 1880 -500
rect 0 -540 1880 -520
rect 1920 -520 1940 -500
rect 3190 -500 3270 -480
rect 3190 -520 3210 -500
rect 1920 -540 3210 -520
rect 3250 -520 3270 -500
rect 3250 -540 7880 -520
rect 0 -560 7880 -540
rect 0 -620 7880 -600
rect 0 -640 1410 -620
rect 1390 -660 1410 -640
rect 1450 -640 3340 -620
rect 1450 -660 1470 -640
rect 1390 -680 1470 -660
rect 3320 -660 3340 -640
rect 3380 -640 7880 -620
rect 3380 -660 3400 -640
rect 3320 -680 3400 -660
rect 1970 -700 2050 -680
rect 1970 -720 1990 -700
rect 0 -740 1990 -720
rect 2030 -720 2050 -700
rect 2460 -700 2540 -680
rect 2460 -720 2480 -700
rect 2030 -740 2480 -720
rect 2520 -720 2540 -700
rect 2520 -740 7880 -720
rect 0 -760 7880 -740
rect 0 -820 7880 -800
rect 0 -840 3940 -820
rect 3920 -860 3940 -840
rect 3980 -840 7880 -820
rect 3980 -860 4000 -840
rect 3920 -880 4000 -860
rect 2530 -900 2610 -880
rect 2530 -920 2550 -900
rect 0 -940 2550 -920
rect 2590 -920 2610 -900
rect 2590 -940 7880 -920
rect 0 -960 7880 -940
rect 0 -1040 7880 -1000
rect 2600 -1100 2680 -1080
rect 2600 -1120 2620 -1100
rect 0 -1140 2620 -1120
rect 2660 -1120 2680 -1100
rect 2660 -1140 7880 -1120
rect 0 -1160 7880 -1140
<< metal1 >>
rect 490 440 530 620
rect 960 440 1000 620
rect 1560 440 1600 620
rect 2160 440 2200 620
rect 2890 440 2930 620
rect 3490 440 3530 620
use nand2  nand2_0
timestamp 1702727979
transform 1 0 190 0 1 30
box -190 -30 350 640
use nand2  nand2_1
timestamp 1702727979
transform 1 0 660 0 1 30
box -190 -30 350 640
use nand3  nand3_0
timestamp 1702743177
transform 1 0 1130 0 1 30
box -190 -30 540 640
use nand3  nand3_1
timestamp 1702743177
transform 1 0 1730 0 1 30
box -190 -30 540 640
use nand3  nand3_2
timestamp 1702743177
transform 1 0 3060 0 1 30
box -190 -30 540 640
use nand3  nand3_3
timestamp 1702743177
transform 1 0 3660 0 1 30
box -190 -30 540 640
use nand3  nand3_4
timestamp 1702743177
transform 1 0 4260 0 1 30
box -190 -30 540 640
use nand4  nand4_0
timestamp 1702729112
transform 1 0 2330 0 1 30
box -190 -30 620 640
<< end >>
