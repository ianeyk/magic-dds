* SPICE3 file created from nand3.ext - technology: sky130A

.subckt nand3 A B Y VP VN C D
X0 VP B Y VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X1 a_290_0# C a_210_0# VN sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.25 as=0.125 ps=1.25 w=1 l=0.15
X2 a_130_0# A VN VN sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.25 as=0.5 ps=3 w=1 l=0.15
X3 VP D Y VP sky130_fd_pr__pfet_01v8 ad=0.5 pd=3 as=0.25 ps=1.5 w=1 l=0.15
X4 Y C VP VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.25 ps=1.5 w=1 l=0.15
X5 Y D a_290_0# VN sky130_fd_pr__nfet_01v8 ad=0.5 pd=3 as=0.125 ps=1.25 w=1 l=0.15
X6 Y A VP VP sky130_fd_pr__pfet_01v8 ad=0.25 pd=1.5 as=0.5 ps=3 w=1 l=0.15
X7 a_210_0# B a_130_0# VN sky130_fd_pr__nfet_01v8 ad=0.125 pd=1.25 as=0.125 ps=1.25 w=1 l=0.15
.ends

