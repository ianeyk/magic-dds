magic
tech sky130A
timestamp 1702791239
<< nwell >>
rect -20 435 200 1675
<< nmos >>
rect 50 0 65 400
rect 115 0 130 400
<< pmos >>
rect 50 455 65 1655
rect 115 455 130 1655
<< ndiff >>
rect 0 385 50 400
rect 0 15 15 385
rect 35 15 50 385
rect 0 0 50 15
rect 65 385 115 400
rect 65 15 80 385
rect 100 15 115 385
rect 65 0 115 15
rect 130 385 180 400
rect 130 15 145 385
rect 165 15 180 385
rect 130 0 180 15
<< pdiff >>
rect 0 1640 50 1655
rect 0 470 15 1640
rect 35 470 50 1640
rect 0 455 50 470
rect 65 1640 115 1655
rect 65 470 80 1640
rect 100 470 115 1640
rect 65 455 115 470
rect 130 1640 180 1655
rect 130 470 145 1640
rect 165 470 180 1640
rect 130 455 180 470
<< ndiffc >>
rect 15 15 35 385
rect 80 15 100 385
rect 145 15 165 385
<< pdiffc >>
rect 15 470 35 1640
rect 80 470 100 1640
rect 145 470 165 1640
<< poly >>
rect 35 1700 75 1710
rect 35 1680 45 1700
rect 65 1680 75 1700
rect 35 1670 75 1680
rect 105 1700 145 1710
rect 105 1680 115 1700
rect 135 1680 145 1700
rect 105 1670 145 1680
rect 50 1655 65 1670
rect 115 1655 130 1670
rect 50 400 65 455
rect 115 400 130 455
rect 50 -15 65 0
rect 115 -15 130 0
<< polycont >>
rect 45 1680 65 1700
rect 115 1680 135 1700
<< locali >>
rect 35 1700 75 1710
rect 35 1680 45 1700
rect 65 1680 75 1700
rect 35 1670 75 1680
rect 105 1700 145 1710
rect 105 1680 115 1700
rect 135 1680 145 1700
rect 105 1670 145 1680
rect 5 1640 45 1650
rect 5 470 15 1640
rect 35 470 45 1640
rect 5 385 45 470
rect 5 15 15 385
rect 35 15 45 385
rect 5 5 45 15
rect 70 1640 110 1650
rect 70 470 80 1640
rect 100 470 110 1640
rect 70 435 110 470
rect 70 415 80 435
rect 100 415 110 435
rect 70 385 110 415
rect 70 15 80 385
rect 100 15 110 385
rect 70 5 110 15
rect 135 1640 175 1650
rect 135 470 145 1640
rect 165 470 175 1640
rect 135 385 175 470
rect 135 15 145 385
rect 165 15 175 385
rect 135 5 175 15
<< viali >>
rect 80 415 100 435
<< metal1 >>
rect 70 435 110 445
rect 70 415 80 435
rect 100 415 110 435
rect 70 405 110 415
<< labels >>
flabel viali 90 425 90 425 5 FreeSans 160 0 0 0 C
port 3 s
flabel locali 55 1710 55 1710 1 FreeSans 160 0 0 0 phi1
port 1 n
flabel locali 125 1710 125 1710 1 FreeSans 160 0 0 0 phi2
port 2 n
<< end >>
