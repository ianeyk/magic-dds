magic
tech sky130A
timestamp 1702726065
<< nwell >>
rect 415 745 555 1225
<< nmos >>
rect 50 0 100 1200
rect 150 0 200 1200
rect 280 1140 380 1155
rect 280 1075 380 1090
rect 280 1010 380 1025
rect 280 815 380 830
rect 260 395 310 695
rect 260 0 310 300
<< pmos >>
rect 435 1140 535 1155
rect 435 1075 535 1090
rect 435 1010 535 1025
rect 435 815 535 830
<< ndiff >>
rect 0 1185 50 1200
rect 0 15 15 1185
rect 35 15 50 1185
rect 0 0 50 15
rect 100 0 150 1200
rect 200 695 250 1200
rect 280 1190 380 1205
rect 280 1170 295 1190
rect 365 1170 380 1190
rect 280 1155 380 1170
rect 280 1090 380 1140
rect 280 1060 380 1075
rect 280 1040 295 1060
rect 365 1040 380 1060
rect 280 1025 380 1040
rect 280 995 380 1010
rect 280 975 295 995
rect 365 975 380 995
rect 280 960 380 975
rect 280 865 380 880
rect 280 845 295 865
rect 365 845 380 865
rect 280 830 380 845
rect 280 800 380 815
rect 280 780 295 800
rect 365 780 380 800
rect 280 765 380 780
rect 200 395 260 695
rect 310 680 360 695
rect 310 410 325 680
rect 345 410 360 680
rect 310 395 360 410
rect 200 300 250 395
rect 200 0 260 300
rect 310 285 360 300
rect 310 15 325 285
rect 345 15 360 285
rect 310 0 360 15
<< pdiff >>
rect 435 1190 535 1205
rect 435 1170 450 1190
rect 520 1170 535 1190
rect 435 1155 535 1170
rect 435 1125 535 1140
rect 435 1105 450 1125
rect 520 1105 535 1125
rect 435 1090 535 1105
rect 435 1060 535 1075
rect 435 1040 450 1060
rect 520 1040 535 1060
rect 435 1025 535 1040
rect 435 995 535 1010
rect 435 975 450 995
rect 520 975 535 995
rect 435 960 535 975
rect 435 865 535 880
rect 435 845 450 865
rect 520 845 535 865
rect 435 830 535 845
rect 435 800 535 815
rect 435 780 450 800
rect 520 780 535 800
rect 435 765 535 780
<< ndiffc >>
rect 15 15 35 1185
rect 295 1170 365 1190
rect 295 1040 365 1060
rect 295 975 365 995
rect 295 845 365 865
rect 295 780 365 800
rect 325 410 345 680
rect 325 15 345 285
<< pdiffc >>
rect 450 1170 520 1190
rect 450 1105 520 1125
rect 450 1040 520 1060
rect 450 975 520 995
rect 450 845 520 865
rect 450 780 520 800
<< psubdiff >>
rect 280 915 380 930
rect 280 895 295 915
rect 365 895 380 915
rect 280 880 380 895
rect 410 715 620 730
rect 410 15 425 715
rect 605 15 620 715
rect 410 0 620 15
<< nsubdiff >>
rect 435 915 535 930
rect 435 895 450 915
rect 520 895 535 915
rect 435 880 535 895
<< psubdiffcont >>
rect 295 895 365 915
rect 425 15 605 715
<< nsubdiffcont >>
rect 450 895 520 915
<< poly >>
rect 50 1200 100 1300
rect 150 1200 200 1300
rect 550 1170 590 1180
rect 550 1155 560 1170
rect 265 1140 280 1155
rect 380 1140 435 1155
rect 535 1150 560 1155
rect 580 1150 590 1170
rect 535 1140 590 1150
rect 265 1075 280 1090
rect 380 1075 435 1090
rect 535 1080 590 1090
rect 535 1075 560 1080
rect 550 1060 560 1075
rect 580 1060 590 1080
rect 550 1050 590 1060
rect 265 1010 280 1025
rect 380 1010 435 1025
rect 535 1015 590 1025
rect 535 1010 560 1015
rect 550 995 560 1010
rect 580 995 590 1015
rect 550 985 590 995
rect 550 845 590 855
rect 550 830 560 845
rect 265 815 280 830
rect 380 815 435 830
rect 535 825 560 830
rect 580 825 590 845
rect 535 815 590 825
rect 260 740 310 750
rect 260 720 275 740
rect 295 720 310 740
rect 260 695 310 720
rect 260 380 310 395
rect 260 345 310 355
rect 260 325 275 345
rect 295 325 310 345
rect 260 300 310 325
rect 50 -15 100 0
rect 150 -15 200 0
rect 260 -15 310 0
<< polycont >>
rect 560 1150 580 1170
rect 560 1060 580 1080
rect 560 995 580 1015
rect 560 825 580 845
rect 275 720 295 740
rect 275 325 295 345
<< locali >>
rect 550 1290 590 1300
rect 550 1280 560 1290
rect 0 1270 560 1280
rect 580 1270 590 1290
rect 0 1260 590 1270
rect 610 1290 650 1300
rect 610 1270 620 1290
rect 640 1270 650 1290
rect 610 1260 650 1270
rect 0 1220 650 1240
rect 5 1185 45 1195
rect 5 15 15 1185
rect 35 15 45 1185
rect 285 1190 375 1200
rect 285 1180 295 1190
rect 245 1170 295 1180
rect 365 1170 375 1190
rect 440 1190 530 1200
rect 440 1180 450 1190
rect 245 1160 375 1170
rect 400 1170 450 1180
rect 520 1170 530 1190
rect 400 1160 530 1170
rect 550 1180 570 1220
rect 550 1170 590 1180
rect 245 1005 265 1160
rect 400 1070 420 1160
rect 550 1150 560 1170
rect 580 1150 590 1170
rect 550 1140 590 1150
rect 440 1125 530 1135
rect 440 1105 450 1125
rect 520 1105 530 1125
rect 440 1095 530 1105
rect 550 1080 590 1090
rect 285 1060 375 1070
rect 285 1040 295 1060
rect 365 1040 375 1060
rect 400 1060 530 1070
rect 400 1050 450 1060
rect 285 1030 375 1040
rect 440 1040 450 1050
rect 520 1040 530 1060
rect 550 1060 560 1080
rect 580 1060 590 1080
rect 550 1050 590 1060
rect 440 1030 530 1040
rect 550 1015 630 1025
rect 245 995 375 1005
rect 245 985 295 995
rect 285 975 295 985
rect 365 985 375 995
rect 440 995 530 1005
rect 440 985 450 995
rect 365 975 450 985
rect 520 975 530 995
rect 550 995 560 1015
rect 580 995 600 1015
rect 620 995 630 1015
rect 550 985 630 995
rect 285 965 530 975
rect 510 945 570 965
rect 285 915 375 925
rect 285 895 295 915
rect 365 895 375 915
rect 285 865 375 895
rect 285 855 295 865
rect 245 845 295 855
rect 365 845 375 865
rect 245 835 375 845
rect 440 915 530 925
rect 440 895 450 915
rect 520 895 530 915
rect 440 865 530 895
rect 440 845 450 865
rect 520 845 530 865
rect 440 835 530 845
rect 550 855 570 945
rect 550 845 590 855
rect 245 750 265 835
rect 550 825 560 845
rect 580 825 590 845
rect 550 815 590 825
rect 285 800 375 810
rect 285 780 295 800
rect 365 790 375 800
rect 440 800 530 810
rect 440 790 450 800
rect 365 780 450 790
rect 520 780 530 800
rect 285 770 530 780
rect 245 740 395 750
rect 245 730 275 740
rect 265 720 275 730
rect 295 730 395 740
rect 295 720 305 730
rect 265 710 305 720
rect 315 680 355 690
rect 315 410 325 680
rect 345 410 355 680
rect 315 400 355 410
rect 375 355 395 730
rect 265 345 395 355
rect 265 325 275 345
rect 295 335 395 345
rect 415 715 615 725
rect 295 325 305 335
rect 265 315 305 325
rect 5 5 45 15
rect 315 285 355 295
rect 315 15 325 285
rect 345 15 355 285
rect 315 5 355 15
rect 415 15 425 715
rect 605 15 615 715
rect 415 5 615 15
<< viali >>
rect 560 1270 580 1290
rect 620 1270 640 1290
rect 15 15 35 1185
rect 450 1105 520 1125
rect 295 1040 365 1060
rect 560 1060 580 1080
rect 600 995 620 1015
rect 295 895 365 915
rect 295 845 365 865
rect 450 895 520 915
rect 450 845 520 865
rect 325 410 345 680
rect 325 15 345 285
rect 425 465 465 715
<< metal1 >>
rect 15 1195 45 1300
rect 5 1185 45 1195
rect 5 15 15 1185
rect 35 15 45 1185
rect 5 5 45 15
rect 15 -15 45 5
rect 170 295 200 1300
rect 385 1255 415 1300
rect 290 1225 415 1255
rect 290 1195 320 1225
rect 445 1195 475 1300
rect 230 1165 320 1195
rect 350 1165 475 1195
rect 230 690 260 1165
rect 350 1135 380 1165
rect 505 1135 535 1300
rect 550 1290 590 1300
rect 550 1270 560 1290
rect 580 1270 590 1290
rect 550 1260 590 1270
rect 610 1290 650 1300
rect 610 1270 620 1290
rect 640 1270 650 1290
rect 610 1260 650 1270
rect 285 1060 380 1135
rect 285 1040 295 1060
rect 365 1040 380 1060
rect 285 915 380 1040
rect 285 895 295 915
rect 365 895 380 915
rect 285 865 380 895
rect 285 845 295 865
rect 365 845 380 865
rect 285 750 380 845
rect 440 1125 535 1135
rect 440 1105 450 1125
rect 520 1105 535 1125
rect 440 915 535 1105
rect 560 1090 575 1260
rect 550 1080 590 1090
rect 550 1060 560 1080
rect 580 1060 590 1080
rect 550 1050 590 1060
rect 440 895 450 915
rect 520 895 535 915
rect 440 865 535 895
rect 440 845 450 865
rect 520 845 535 865
rect 440 835 535 845
rect 285 720 475 750
rect 415 715 475 720
rect 230 680 355 690
rect 230 660 325 680
rect 310 410 325 660
rect 345 430 355 680
rect 415 465 425 715
rect 465 465 475 715
rect 415 460 475 465
rect 345 410 415 430
rect 310 400 415 410
rect 170 285 355 295
rect 170 265 325 285
rect 170 -15 200 265
rect 315 15 325 265
rect 345 15 355 285
rect 315 5 355 15
rect 385 -15 415 400
rect 445 -15 475 460
rect 505 -15 535 835
rect 560 -15 575 1050
rect 610 1025 625 1260
rect 590 1015 630 1025
rect 590 995 600 1015
rect 620 995 630 1015
rect 590 985 630 995
<< labels >>
flabel metal1 185 1300 185 1300 1 FreeSans 240 0 0 0 I1
port 1 n
flabel metal1 400 1300 400 1300 1 FreeSans 240 0 0 0 I2
port 2 n
flabel poly 75 1300 75 1300 1 FreeSans 240 0 0 0 Vbn
port 3 n
flabel poly 175 1300 175 1300 1 FreeSans 240 0 0 -400 Vcn
port 4 n
flabel metal1 570 1300 570 1300 1 FreeSans 240 0 0 0 Vx
port 5 n
flabel metal1 650 1280 650 1280 3 FreeSans 240 0 0 0 Vx1
port 6 e
flabel locali 0 1230 0 1230 7 FreeSans 240 0 0 0 Vy
port 7 w
flabel metal1 520 1300 520 1300 1 FreeSans 240 0 0 0 VP
port 8 n
flabel metal1 460 1300 460 1300 1 FreeSans 240 0 0 0 VN
port 9 n
flabel metal1 30 1300 30 1300 1 FreeSans 240 0 0 -400 VN2
port 10 n
<< end >>
